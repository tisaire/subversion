��/  �Xt�`$�����My<~}�A��5@%z7�FH\�0��-�9EMx*1�s���v�G���n~����1cg�&Ft��ͽثc��N�i\r���y���AKK^�z��U��Z:�;��KP�B ��N��A�[� ��P4Xi�%�T��x�Y�c���ۣŤ�LV�laD=tp8F�=�}A1��=1�<��xr7�n�?��;�MHc ��c��Ɨc�ɍ|�w1�ag�j�J�gDBʚ��n�N���a�� Zs��Gb��'�[����_��.#�2��*���|�PNž�0t��'�֩�X~!���i0��A��-�xI'O:1�T���v��W�r�� u���ڍ3�����G����Lֿ�^PQě��zg�nJ����*��EV�I�����u�杇�e,[��l��9Љ�`u6���4�
R�ox�uT\)F�^a�¦/��`ɁK�<��]Ñ�tt�GGe��[�]GO���Ŵ_Kb��f�Ok�i�(���\�,��br;ғD����1�Q������$7�N�����S?L��:�sJ}��%oy��������3�ڴ`��?�le�9��<m�P�y�!�!��sN�E��k�+h�602y�n�AtW�����V��N�"{�042'3����L��l�d���E�3�����Li�&3�����o�����Kk��:h�A�,:qoB�qU�g/�_a1hl���vo�$v����3��4�?-N[����w ���nG2ڻfod�<m�)�������h�x���n.��q��R��^�w5��76�� �8�m<�.U�@�:���i���jH��Ex�Ю���N����.�5p�V�l^�������Ft=֧@{�k;Ee�y�դ��K��Y%��b�ĸA;�QC:��������F��c�A��д�~I��O�,kL�S���q�eH�R����܅�g�2ۺW�M���?�!���;��b��\v|�d����^^�Ȱ�[��r;�e�WN��b���t�w���KĬ��O�y���-�gYդ����m�3�Fbպ����u�@�TE����Ȳ��#���I�>Dں�GgQ�`(��	� `������H�p���X��X��i9p�s��jCLa�'rg�_���ZǪ@��fͨ-�����Ia�a�i[�73����$��.�5��Y�׼2��KÒ�y����$��\�M�/�s��s��4�37��Q�%z�O;h�T_c,�uL����I�<�D] �L���Y�`~'&)��Yb
�����%�ㅲ���0G�wUۙ6b`f�_!.:("K��Z�=1�'T �p,Q3�1�/���b���fī��ײZ\�m��B��s?��:v؛��ގ<���ޟ�3i'�a9
������l�5=�A����;,¨����ۏCC��}��P~
�F�ݔ+�].5��-AJh�]6�����0	�~�2�U�*���Jc�K��&�4*��@'�U˄YΩ�)_�}�˶Q�� ��5��6�:�?���B����U¥u���?�Ҭ=�>�V!�Ã��� ���S�4���O2�A��.��8��P=�V�8	����i쥟�;������_�B]�@
���23��`���6��'R��2=�껟M\{b}7Й����֕����!� :��Xh�`��)�:Y|��B��b��#JDG�kgjꅶ9Q�+���������������f����x5���wK�U�[/��xuv�t�((��]2d�;˶�O�$&w{UQ�%>���\#!5�*�LI?]c����^����?�s�^���Zf���Mw��"�WSP`�9�g�nۢyXT�g֬�-�i#��h��ʿ�py�ِIP�q`�����8}��h	�(�ei@�,L �ҽE����~{K��fj�E
��T~�T�nl҃�&�W:�/�j�mIݡ�
����P��k%���DN����-�>��42��G���9yZn�O�祗)"�r;�s��O41�>O�FAo�ߗ��3=�Pf �e0�l	ca4"|ʪ�^���/tUw�%�.?��b��Q�ܷr|P<��@f�8���Ww�$�^�A�g9�it`��<����k���P؞d��ݝ��gS���ۙ1�^�U`��j�x�+�1�◩}b��ဟ-Ƞ��q
����U�p�CʄȄ-�Li��,6�����2D9�3�+���X{��+!	��|�t��g�<��8�@� ��"#Ь}�^��n�M��$�]㴎8�ꬠ��l����̥|��k�BF�c�!��z�L�9r��a��]t/X{"�(�9��ww����h}#Ty9�bi���J��k�qO�(��}�*[�}��^���^����5��i�` T�#��Α�Qۓ;�<�W������s��U>n��˫��WFF1��FA�7F��y�%�pu���톖_��2�_�n2j2w����߲L��o�P�!Z�����霾Y���vB1M�����=�>T�-]ݦ/��=�n$g2�ܥ�j�O$@�VW+��ܬ���Ï��ٺ�+@d��}�l�$��K����#+��h���xW/�����;����������
�}=����&���\��R�?�i��HS�ԍ>L+�8�d����_���6wt���ZՋ ���铫���|&|��ʂs ����\����!�~GX�/	��G�J�f飝�L�э�����Pߛ)���:&:�|L���u��Gd^��l�����|2�
�al@�u��iw���O�>r� AS�^ ]������~a	gA�B� �%2�������J:ͥ���я�Ws����~��K�^[���Y�����<5�� C���F�Ƣ�C۔^fwb�����2�P��֙e����F��a@�(Ⴇf�;�6~��v�0�bYl�g����B/���=����0����&���R�Y�]�F����X�#j���|7����_�j��B�o�s�[A�f#��*�o��Ck~��j:X�_o�ao���4a\�+]����K��M���H��&�k��?~{jµr�2��%)#Y���&{�ivp�bG~�L��b�VQ^B��
���;y��.U���3Қ�����%�2r�K�{U�7���qR���\�k9[ž ���/���i���-ѕ��L��V�^J��u!{I'1CQv��@���'�e��<�A涏�~п����:�uK
���	iv�R�!�-�1p�ߎ�3��'�i2���_Z�,���(��'V\�?M$�.�@�TtNu�v���ӜW]W΅�N2qA��ۥ8����h.8l��2�9Q#��sU=I���K�����R�` Y�=�:���<��@�!6e��B7!�I�Z}Yڒ<�O�u�D��?|ϔ�1��HƇ-!��x�8��Y�K���A՘5����Qsw2*�ߐ��X�/�j	���� ��=8t��js(��e�V��XM����l��F������t<���^K�Ą���kJ5!_��XZ��1 a<٠}��2A���	ȩ�hZ�����v�V�0���ˋ��>:�+�<���A�6^3�r�'8�6y���$z��%k����O��cGȗ�<~���Α�įD)�H����+|�v��AX�ǩ=<��௨�x!�����b
8������y��Zߙ�����FM��r�Nhw��J�:�>��N��=־Q�0?@��i�9R@��u�>ؤ�U%vJD���s����J�'T{�:
��E$x7�K7$eq)��u�e�vRV/9O��ݠ!���w ����\�x!z�v�+-�atҋ<p�;���v���0�w��{	O~q^�����K��Y���ua'$�X���Z�w��Vk ]�l��<�}I����F�ͼf�#hg��[P�5]�/�5��3׼�$��݇��5���ni�����i-��5-��IE���QxI��s�o��rž[�g|�~��h^v��6u*��F�}��b�Qش�
��Z#�=��s����[-C�8�1��,5�4{~�/��|>\��X�����o�a�m�Z��t^�/Z9a�Ss���ΩAb!���Q�&�7�8fS��U�=%z(�n�o0�j&^h�J�|�O)����0���T���<.hM'�,�Z�ᔸ��q��ﲑw���n�E�.��C���V�:t0���,�~D�x5�]�����Y���p_����p�.wW�JO��u��-g��Yg5�\��C������J+nC�=�t�I�~z�%�P�'����ۭ��靵��C�/.l�0���>�n=X��**��s����1�Wk|ddQ�\`�r���CM&�s��w�ǿ�C`o+DJ0ٝ����-�J��ո�M�������&&'<3��S�2�1�����L���yH@�%��	��V:���޲�i���!����YJ�:\�9qrO%�i��E�x�_�Y���k�f[~S���h*"���tk�T.g��T5=.I�����
�D중��c"O�G���Gn��y���-�-s���"3t�pq��ԩ��#ZF��T�d0��nt_�JQt�M����@��ԚI�Q��9r��Q�ߌ��y�>>���X���C�h�`�v<�k��*_�rl�O���ޭ��*��\YjR}t4��O����]��賿8r���
Cl5q%�=ޘMŮT*��>4�Z���&�)Jv���K��g=&��»���zr�d�mZEX��3m����(!Co�u�=�� ~��#5�l��&o��'��}r5�)�*��7����J+���C��q�k��!�r^Wύ��E �%a��NzT�is��G\g���\��p�S�~��VzO��q���N�-a��C�?U�;2���`�0��=!Ov|q.��D�@��!PXN#B�<٠q[��1:f(�����"�v`�Q��ɵ����,�2�����| ���c�hEڵ��uJ�֙����M ��9�j�\n
�����~x�1@�0<fJ�Ӯ�r��ױ;`�D#�����1�$R�B��>�i�v��ڣ�k�ǿ~�F��N	�[�K����Ce����knuޑ�?qAX�=���czi�0�%f�K����<����o�,M���^9���ΡFb;�s�h�H��W��p_�w�Ћ�3̭��y����YUj�q�9zSW֢�	:�-�Rc9L���(����W��8�E	J޴Ґ��{�h����F���ܺpH�W�d.x�&=��L�yg��W���)�C��N������M�[f=�_�FZ =���r�6��� ��acD7ØeP����re�gbDhpZR�|�h䥠ϳ�!���K�b��Cm���4�K��A���M�Y�X��l��tD�i�mAR�]0� �w�]�����Dj�?��\�c�v<�IL��!u.��ƞ:��
�]��S�㼤�v�\�t� ��U�	��cjLe�,~�)h��^+�����ow�Y�,�o���d�.®�o�10{u�Q�R�k�h�%'_�m �����(
j�Ϯy�"$v܉�7oz�<B��v���T<�s�G�&��p�ʻЮ�l�9�'�'Gf�nw�eAq�	��vh��@��vG�-q�A�Z���{�d1N���!j6�75l8���i��+���V(���?{b^���a(W�nE6��2�a�TZ�/=?%:/�@Ō:x��:��p��>����9�;;��T$���{�;vd����n�x�&{b
#�l��C��� �%�p��_zeZ�ƍU5E3Z�A��;�U�(�xv	�l�4���3��hޤ�TD���{l_%t�O���&9�`>�9�ږP%µޘ�"*��r�O��9o��Vc>~�����12Q��hnE@;y"�gyt�F�ۅ���o=l���l*�-�x������T}8S���+���=�6H�)R�A穩ˁ�u`^3j�t��9u�$#���@M�W\Y��پ�1WM�d2�ȗ-Lspa	�������'�'3l-�k��]�T������q�.F�0v�P=�oGqF��@�]�DP��b�#u$nW�1lsbM뱑�xFM�E�8������
�0dPu8�X�*+�ɡ�`���:u�?C�䑕���s�K���x���gŨa�zYD�3g�#x�m�o��L�2=�ds:= �����utO(��\'���Ox�̺��9#�z98 pYpz�?�73���5ץ�elgt��v[n~aW��t�1�n�%�P�J6�b�d�� �%q���PJT��#Ա�u�@�R�Ȯ�sMO��"��;Br�fk&8�6��-|����|%�����cj.�\ΏN�C�=��`��r	�����"�L��#�.��D��`�6�ƒV��CIh�~;���Ξа�R$Å����'�:% �j�a��_۲���	h��Ś�w2g�9!N��8�QF$$�z>�҅�d޹�b(��C�'���(�voyC���m@q�HE��"����f'�q	h%^\�n�.~/��]`��}��Y�w�(�[X�M���,E�,6�u�d�ͯ����HM�K�T����t�!�u�h�!�}?XcG,����z�Y�L.[�@��O��w�#LEX��<f<}cs�y�_����h8�{�n�u&���*��h��ԛ�+d�{͟���6@� �S���roI�D<c���՘1no2��{����q[��_^wL�Ə�<W�������N7P�n��#�'�>4�7/�/�{�'�'y�;ɩ�9BG�zU���i����|��DK1�%2S�|yVp�r]�ɠ��Ƹ~sH)�@��,�qhfշ���u�f�1�N���:�'�Q5s^͹�-,�~����%�RcQ��.}u�w���]��9��|JT�m�
����o�7zѮ�)��졡y럀���'��tQ�w�/�@�8r�������r!H�j��*<�h�踱��P�q ��C�/a�#M�E��ʴe�L֨�Y.��/H4Vph"���s���/D�F���#���:�8�ɀs�In��L����,� 3���Le^|n7�XѺ�d�}U��:���ɐ�
BT�_�#'~\1T���T�l7���&���(���a�>�;��T�Z�.��	���ӫW��.��(x�)[V�����b i�1�)�!F�g��;��H�4h��U8O�K�e3��&߂�Ků�xhީ�`C8�!�Ǽ��j/`��4��VK��k�o
���L��.9^ڝJA�Er���T)$̱��`�Ȭ���߭ӥ��1�OORt���^�,fG(oG���XS�V��=L&�~v�'����ܞ%�S4�gD������o��n�y�l,��l�}�.#�'Byfb9,���!4�6Q�����6Bݪ_�{����ߑ�tNp�xVOj��
�lA8����cW�W��0�+�3wG��)�i��cx˪�r HY,��$kǓ,Ĝ��U��u���N���R�	��	y��n��;���бuc��Qp>�o�r� ��0ꐲq���H2.S91��gu.�'y+��N�B(�(��V��*~���v�{x|��h��+-��� �&������u0C �]�L��5n���!���z|�6��5��s}�-���\��І+!ݪ�B6cVŨ��lBؕ�'��SP�i�;�����o�N��KfsR�:�}��j-@(!�!��g�L��9x�~�����n���&���RƝ�TY�6
'����1L��`�2Ld�B���אEN;�X��#��8��Z1r.�N�Mt��^�9n���gJ�:Ms�~���b����]�u]��-�̪�=]Rn[�-�h���Č��WjqE?C}
�C�n�Г2��?ĕ���5˴�H"��,F݀QA��B�����!�pH�'&����r��c�Mݸ%�ܧ�<��Kuqx�X�àΣvm�1&�9�&vʣ�,��k��E��`�i\�6[� IE1a>�B���N��!�.2t���4��H�S}x��q��Q��ق1Q��F{��eD�Ϝ����� ��@���#1�<��½ �b��*�%/��e��e�sf���2wurR��,_���LUIw�۠�	� �=��k�}����9�_c�����;'h]�mQN�f�����L�f���J�6G<Ҷ{�>Kdٶ�F5���f@r�N��)�nUq�����cbǰ6��#��K��줃=Ã9}�K���c'�Q��}�)���f#�7���=Ӄ�+�7�j�`�}y��$
��̃�)��h������Pv畼)������	N���S��4�a�mi)�m��!Js��a4rϷ3�v�u\@Oyisv"0I���-R�l���EZEs��ϓB�q뎝|��D�c�;Q}�������=��i��Y(�X!����R��y���ǍP��#3�Upk�,ꝝ؆
"�=�^K����l�z��Q<Ʀ~�+���2	H�A� �s�����p�����A1�Y�@���JL�X��6-�[�O�`_��j�o�B�I��s�Ɏ[� ������4��Fj=�KR����&�z��fV���1D��{�h�8h�jE?Z	�U8|Em�}�9�Ն���,��Ք��F�a���l���N���[���z����N�S­v���EʤR?�7��M^%����z!LB� ��墨&)�5�G�:�p�;��t�f�5 ��*^�������Sv}��/�=ޕ�������-��z��pK��c��K������$�(���e�Ev��q�@��6���5�k<��o��*�'u��ÊvI��R(9�6OE�������@�3sQ��z��e�^�1�O,��+�I�ų��Bvx4�zP��6q!y7^?�]��m�,ic� ��Q��`@l�eg��J�n�}�Ξ�������!�a�o����P�^�)��*�6�H2Q�h����h0\`X���ā�ޔd�I���M�ߒk�V^?��>߶�?ͯ|^�?��+
��R��4�S�Mp&��'8�� I~�l.�J��7�^�
�0M��=涸 At�Bu¨n����>j+����ëM�J�.��1;� �D���(��w2i�S��;�
�:0�-�甗$a~���c�$�g���Oi�ᄬH��*��o$h2)���U���g �K�ʌw�����P�;�F����۝I� �$�#�Є��2�}<eGJ$����ؼ����̧��"�
�7ˆH��~=u��@�k*�g�HҖV�n�`1�z�e��#�f0u��O�_�Sa�Ds�
�w"38^�����;o(%K�]�W�9��������R9�F����]q�7Iֺ�%��
�^o���p*������.��օ�������Ǒ�ȚG��8_���N�ߕe�B�1W#�4o�ǔ@]�D���Eo�o!�0�&��w<\�H:|t_<?T���*�U�D	Na�"Ϯ��&�?����S�r�V�tO�O�k�tu�n�o5G��Ao�$`+��嫋̷�E�W>���t@y���L�fwy���Z9��U�Z�l'/�N���l�9�<$�ʘ&�H�P��f�h�P��_Y��æ�kU1������uY&��c��G���!�	D�+� �H�+U"*Ջ���çTg�<)��7twp�b�pg ^�Jݮ�a:�� ش�!�����0\����0���C/b�!J��F*��ѵt�ۃVjNX�R�P��֭7I�OX�gՐX.�������0�^⒩(n�0_h���DeBT/1A��Qa,��U�J����ru�S�)�i��1��#��ւ+��j�ڇ�3޶���fW��|陋l���-ko	RU�\+��ԛ��F隂��(��V�
��4����Y�ID?
�����L�3����B��9:ʦ�����Y���1VHtq//��fĂ�E�4!62��ׅc�%q,��N�X�\�l#e�4��f����rV�G�)f2�:hdgo�`Qܤ�|6� ��+�B_��Y�N���87K�5F�����D>�U�2����4sǵ�{얡�6����*W1x_��Il}͕����:Ax��W�ܷe7
��+<Q�h0i��<ɻ�s�xw�t�RIw�6��#�ʮז|�#�8m��a�Q٠9N ��{zIv���m��}2G(;��'S5�`��15�Y�#�u���j��%�h�mVS��6gh]Dр�4m]7mݭ~�hQ�	t�����U�p�%6\�(�.�H�{�=�{Y��W��f*����m?81�@�;.�vrJ��	틋A'_�.�}]ƴ#o�TrC~�	r�����A��Z�����.u)3QP�gq��.~f_���K)\�P�EV�󖇇��*�~��L���_z�y�j��z��T�;1ae�U5��x���\,t߹������	���Z�{X�[
�>X����������"�3���G�9�)��-�B"S����m�
�F�|�����t���Ȃ1��Žφ( KFk$�0�b6��[�1�Fv[0���,
���#Ri��O���R��v��	1��8�O�'$X0�1����&�\$��q�G`=��\*����5�&��̙���X��Z�W�~��AT�>��p�Q���?@�|^��U�#�u���1�ɫ�![Qe]G0�'��0b]�5�E9�,K������Nw4�D�~dÇaՀ�Z�(�w�&Y>�J�
�#�&��p�OZi �����"ء�]�i�����k*AOl@=���{�ٟ��%�Gx��6�s�����9�����{%r�q�ʏy�&ѓ��gݗ|�䫸׶�F���}��3h��mDnw��E��f�*e��P�\��G��b��˕HΪNF������9>L���]��N�v�Y�s�!�r�W�g�s�Gп�_y�M��Һ}Zi�Yo<q*Y��}4+8b9}eŻ�"jc�s
��M� ��l\J�����bE�T�˴�*eD��/�~��[R�p�M:�$�� Sݤ�t�k���&Q=�r[��=)Xp2?�8��k���WD��}�꽃�m�
����o5=���R��;��};��x���#����y�lŅ{j(/�B[$AƧ�N�f:yvtۚ������IUO�T��f�(���$>�o��!f�qZ���Z���������W6
.�	-�F׏n�X���J�]t��J/��Li�;Y���p�WY:����H�|thb�Y\��8�]	5?�Hi���$!�9i�)W��T1�KL��%���Q�p@.�C��	�&'=E�������qٿn%Ƹ-��ɉ)yJ��ø����L�L�Ń�rTn���̀�xZ�H(��ơ�c?k�)�S��:�����G��П�+�LD�װ]SBFC���`O������`�ȱ4��l�7qn�mY"v��������H����JP7�D�9��2ڸfaf�i�z�wjأk�ԏ��>�k"���"5���6>_o�|�3L8<��[9�#<�WA[Uv�>��T�ẇ����L��*G?���9�Ac�qd�k�Ɲ��x��q�
�����:��q4������Zk�d�\�ؠĤ�x�*њ#��J���xdIͥ7��%��-՛O�"��X�W6��n��2�s-�~A�L�8�͜��2w���DGC.�G�m�W�T�v(=w����ؙf���u��lՙ$a'Y&�S�}�S��)��e����ʔ��e>W���E����D�5��|����mC��C�=�)�QoV5��6��՘�����Q �Xp��ߦ�-d@׵��kOv�>r�Qz	�(i1�H��G)�&4��M*TqM1�w3^� bX��;�Kg�[�/�ѽ�29�_����>��39���u����a��ȏ2!��:$���+��J��ffb'�M6�Ɯe�=	1�l_/@�"����n��~[ ���d{��n�ާ|�̷t~����/X�i���w�̰+�*K�5��͵�t�Ur	{����I4��Og�@?/��i%�w������%Y�:E#��_�LI�6ȉa3�QL��ɻ����}	��!`pmǽ��b�5R)���z{ۮ�@i��D�9	�%�ڌ��I|�cXs�.�ӐW���y��z^������;C�����������(�a��]$}#���\���Xb偩�iE�gx�Օ�!`�^y���$fX{4��9�D�<\KO(�r{_�)d\�a}��v�v�A�8A�9)F�12ᓣ����_yc}�f��N�H�;2.��/���VevB���47�����l���Y�u%��	��L��n�&��6�LS#����vw ��k��f]5�2�u����_�Q�4� :�`+�v��qo��d9}a+���|��nc�[4��u-�/�+Huh���I�E�E�u:�n'_f�M�����im���C�,?�jo|���L�j�����ǐ�.<ӯ[�C���� _zY�S�H״E�:h\�#��<U)�J�L��2Q��5MLv�*GɆ��\i�kh��7[J�7W�yʱ �+���U��	��F����~S�>,��"~v/�UN��%7��K�K����CW�˅�
ӂes
����Iȿ���g���T����������L��M��=��#1�D�$�+S��]��NC*���r1���P�1�n,��-�RP�zϠP�s«�f�OGa�m�B�d�<p
Ք��	)�29S�2��v/ϡI��}�R{���l�P�<,q��υ��q� �S�/*Js{�8n:���ߋj��pi�6�L��!�����b���-�*���{����SN&u�d2��0�t����~�^ɜ�G��a�Q��'mX^�l��T`�O�����?����+���F���?�}���(�Ա����s�����c��J\��)O�]&/K��eo&�D��~\ӿ�o+�'���-�4H&�fK=la��y��>�I��9��/�2K?y��[�#Q��n��s�a>dGEeI�.1��~F�����~U�pe#�C���-��B�œ"����9�l`<X��[(�P��� ��?�jP���槆����:���Vpv.rъ0�`z��UD�D�mH�"��Vw饬��˼��n^�dꍝ#��*X⯧z{y�w���.��c:�W�c:?#����t�����Y=e��Z�����=Ob���"�(њs�n�_	��9�S���3�R�b�����h���&v�4QKm�.nڟ7�rZ��N�h�!yi8��+M�H������qݡ���
��i�*�9t\��`'�ɼ8�ģǤ�u_{g��A�`��E��n%�Ό�TAHب۵�FL�N]�±S�J[���a|�����w�|��?�N�u�Н?�&��������O��� #}�}��9�c�UZZ�sL=���3N;���J5���F�B�,��	R�@F��W ꨋ0r5ޏROB#B��5�)(&[�(�!X��;��r!d�L-�P��6i����t+�.��
Ȉ�b/�Ey C,�{.�7nT:��YU}@��2������ke%;h���/OA/����Ռ��Or��V5r�!���{4�_'Z�fY9cjǋ��㓺wIF��7�E��6O�1��T����%cG�$ҫ��FF����|���D!.�ו���p���1�SE�ob�O9a�5�V_�d�� �~�[�U$�2�v�*�2ے%ˆ�y�39�r���46?i˹�.i�k�O�� y��)�.�8����Oh����q)E�������xWԌn����nM����/����v��G�"���u���@8���Gj1��{����J]4,�i4M�(��GjU�qְ*��1�� ���{Rt@I�;K�|fW�b��*}�� ]��;�%X?i��n�$����{���B���)n���Qd@����+zA5�g�hJD��T�Mr�y�=-�g��g9hG��d���l� �p񡈼�00�/�b�lp`���s�f��c�o����
����k��˂�7==��Λ�=Y��?lD]�mwV���_"x�r����tC��&K&ou�O��o1�U�k�����T/C�R� �2��zgg�)���b1�`�oQs˹l(�+�����=�		3D<^h�@8AE�M[r.������Z>�C��)�}e��Ǖ�}�~���8D�V�"/���5u'�Mܩ���v�\B!�����T��o^�JS�*x��U)k��!R��nzbz�M2;�q��閁���y<���L�:���s9�c�l:DZ�5�h�����xL-歳j}�۽cq�N/�s�s��R��v�d���S�/:�hH��r��Rks~�;ws������8L�n��a$gȩ����(����[�]8Dd�qI�vV�k��-��
_��N]���v��c�ǁb$���+Ľ�6�{�����������u���)B��2㞒��(���T�&]I1(*!�N@�7U5x���ץ{��c��������&t}9@�ԗ�b3��g�i%������(|� �:�gKtDӶ� �- [�j����2�%���7�H�{�-�
X�k>���c��S���$���_�BH`�'��IA[�f����t�����`�9i=������c��T>&ޤ����,h�o�7������8P�mT����]�D��8��~Ķ�n4s��P$|J��6 J��;�3hd2��9s9�������7�������ɬl\T> �m����biDob��G1tW6-t�]���C���}�*
  ���}�h�ؤ *5gM��:���(U�+�\4��"���E�r�����j���'վ�;̅�_��!Im�B���1D�;�-5g��k@ք��L"��h��oc��R�˃]�终:|X�z������xm{xr˼���#���K�(8�/�}#l�9s����5N��s�&���r��=��T&���\�v�3>;��-VBWrd�a�j��Q���a
�]̲��O��@nQ���D+��!ڞX�T�8�s�ұ�Btݤ��``2�܁�����.��N!�x7n~�b�cx�o�肈wF�qV� �L�~-LS M
mB���nHh��#�5�jV5i~;�4_7r�|��EG��ash5X0��2���Is�h�#Ռy����s���n����a�����aEuO ���mu�'@���0v?h8�z��T
D{��fȒx�t�j:�Rk�g��������|��t�㬀�gi*X>4"֒Ӯ����`Z�Fd#,׽�P~~��E������������6P�t�z�a�
�0~�MD?��͕�{84���Z����<yA�p����M�㐖�ޤ;4̩2,�LY�[�z�>��7L�A}]H*@�s�<�Z,��*Ρ �ޟ���u�A��u��H�R��jG����3x�ٺ���8{������i�twt3�B�/�Y�uK�*d�����@%w򃱨-a�g���[0�ͳ@�	x}*ܱ�7�@U�B�_ό	������&��_�6_dId�EVD [@�'#��s@�ۍ����K����NȜǚ�>ȘT��VB/u�\# >�·�4�$�q5�)��<q`
<d4J6�˂�80�6���z��5��	9���#�q��v��*��w"������g��~7��٠ET��OqW�*Z1_�5�����|����������Wf��5�)�%�k���υ����G����{�ݺ�>�"�6t.���1s�e�+_������Z��m/��i�d�/K60о��q�2��藵��\�Pn�AQPV�$5���u�+'$���t{�����yԭ�Cn�*�3�a�i���CX�'#Nu��lM�tJ΂ �I5���
���E����QT/���S��DN�K���p v���/�#7d:��C7gMQ���83ڄ�? ��*x�Mi6yך��gY�9��[��-g�)���F�t���K6�*C[���j=#G�hHL�Z+Z���c.2��΂gя�K��ɽgr�T�0�+�J�N�;��Tz'��m[�Xy`am�`��r��į	1���g�{����3.�5���a>*$����W�Ѻ��4��l�{��-�x��*�DB�m,-X�g��~[��W�kn'��#��$��\4v������m��F[��B>ѥ��a��1��d�"��GmLȶ7ҵ��@X��N+�Ǽ5�x�����B��0ht7�ˤ#[fZ����1�6/5��K�p���o,^�Cm '�vkĞ�B��N�
�/ٱ�yq�s��&]���i��u#{Agx���B�m�H����T2��V���-�0D��Z5��.��E��-�:��˦1�¿��;��]�s_	�u(�R�\L���ll����I�١Yʵ]�	����4)-�<�Hm���,GeV�ǐq >qz|.?}d��*l�S�v����;�뢿�����96�-'�������	�� �Z�D��Iwr5�n���,w�$�0��uN�����5�81�6�"���G�GcU֣�j]�tӸ���w;�<�ok��
`��&�pp1���"��!����8�j��(x���kP������]�����S��e�&2L�s*B�)4�ُ���{R6��+/�9��Yߪ���y�Qn�,� �c�^Sv��}�v��TC[<��VΉ2�@�X+��ы�N��`���!]bA�&ٟ�=��l#�FѶ�Z\�dx�;��{�F�D�ޘE��w5��o��� ]�ΪSW���Z��6�	H1��W����U���:������M���Ry�O��V6�m��0��ۜ�ޠj"��Զ�3�����3�8u�L�̓Q�;'��K��G%���mK�զ %JMʽ@&^��㓅)��P�Ӿsu��b��Y��{Yk* hP�{�N��WT��|�u0��)����Qط�b�=�	��!��vA 匥�
��~���=��r����](͕�`:r��W��.�H�7ւ�q!�ync���H��������Ǔ�	O���׺�E;k��Mz�7'N��PK��gu�B8�j{���kJ��a(!4�@���j���W���ꁧ��эE%n��Y~��R�,۸���؁�*`J�C a������4��t����ƾ��{Z[탾n{�	�9��!Z��t��͈�[Utש�$�_��)Of��A�vo��=k�u
1~n�A�7]���u��Z�2Y�y��nZ�8Z61����N�Au���)&�'�l��%O�(y��
�7����e��C,@ڎ�G����_)3��j������v�V�	2^I��H)��jS�:��!��]��ۊ��W΍���ܕ�d�H�WE02��(��M��}����h�ܣ������ƿ�>m)���@��f�����f�vVv~�e<�?��Ӡ���ݗq�'�X���B�l�����@[��z-�
?��H��������`�yaK��d�rj� l���D�$/���mT������	��@j���W�s����ۋ�^� ����fT.%���j��L�Y���$�����)��lVI�g^��XM��]*�����U`���&����_CX^|Kȏ0�w�mPY<�DHA�C![��͈��c�:�M�'��`+�a�ٳH5~V@���v��5!ݬ�d�Ɗ�A��.,Հ�5��K�xiOlC�'��w�����GC�fQH:e^س����λ��C�����M����\�u"Yw�,�0�QL�(.͋�j@�i8B!&=�����3�b��7�O�|�C<�|����Y�ZO��+��s�@��d�=��3���0|�_%Ť9�ݱ��`}KB�2o��^�+��H�R���b�y�nu�ne�p�j?���@-1�{f��א��f��QY�Uڂ%�3Q�]���
�m�Q�M��U	O-����k�A��R��u�ٙcWŧ=�@�P�Ά���fo�?��u����0*%P��-�;�m�+�#y�рo�\[4	�ԡ.�5!�Ϳ�*�cFX�D.���问�@(ޟ�N�M���(�+®@�����)�M���J���Dq��-�Q�F��=)����S����q�G�w`�e�C�!����NW�OuۛU�x;d,���f���5mV���A��@�6;j���E�ƪ�d�O:��0fX����� j����?����?"R'�}m��������r�о�.mY>u���G˧m�H�����@��F�(t��!1tIcHy����>bL�ٛ�>1��?�����3�i���++�f�CV9�(�fc�L ��J��b�RdD�cd� �!�(:h��Ě0�JH��=�Gl��u�c�����SJ;z�X������rj���>����T��P�6ż��/R���4^�<�bO��k�:�O��wJқD�K�>
{�P�e�0���^�[�����T���S�_�ycGt�|�GXD�
��iY�|g�^ Z�x�|��f|oU_�4L��/j����K��X�Ֆ�8�xՂ��ڜ���i���������d�k�įsD���<9��)�l�k��Ȃ�þHY�{��on�00�u�����_N%]moW��`P�4��q�Dm�� �OO8���~e^ɜzb�Sc��^z+����S>\)��£��l������� ڙ�y���N�^ۀ~����LZ|�����M��MV�Q1�Ȉp�r�4h����V
�G���Ƞ�k��Mien[|�4�>��!��
�-P^� -[2\����IkGy�ӹ��Hqs��H���c�� r�} �O]"u��u������$0�[zd�}肜\�+xa������0���?�T�C���<������}��ɖw��#�0!I˺��8� �F�j�i
E �|#*C� �ԭ$�W0��z�M.�/9������'B.q&�0��OU���U��y)�3���V���d�$L�z�30X���B`v�T��Wg3�ه'_u�<���CS>Zӯo�t�4&^���\�H<$����tE�������_�t*Um�FN����?�[�)]���`t��=��c��k���8�3li��N���/T����R�;G���i��\���%����]1Qk�����nV^��A�K�L|+\���H��N9a����]=wv�[ȴ
����6t(�-�Y��$v�z�I�DV���g����I�N1�����o��/��.7�3�隳����",/D�GOʦ��ཱུ��x�۶1��
�D�����H��ix|ʵ��������[���~b�h��8i�p���@
��+4:%�oA(�2\��va�x�*u-+�|m|�|Ĵ�n'(��WU����@�O��8!��*Sw}E(&�IL�{:�\�d.��	�4qP��t	ra31x�����l���_͊w�dh�����ڕ��Q�O,�D6�V��/Z�'n-���H|n4�lb��5��z�/�rX�c%�p;q���e��=k��O9���p_8f)�Yg �pHe���{	s4�%Y��\zC�8e��~mܨr�%YQ�K.���w��C�TH��*��[����� �- {��<�ƺ�N�
O#<����6p	���3��&ߔ�	���-	BT��7(;o��u�&���`�߻)+䀕�	�j��G������EVإ(B[X�� Ӏt���I�����I��7#�Eۦ
TFФV�Am�O��{w��}gDS�o/��A���b���r>i����=����'73�j��їjRl/y�y��,��v���
��V��}��c)�N����Q�^�x�bg�nH2׳vwQ$Xl��*�h�_�d���G����/o�C��?��M�}�V�M��*�yR�����l��5��.��؛pƌ�۳-��yo��szo!�p�-Iߩ�nY�ֵY٥��� M���?s¢��ԆwL8��o�$�`�-�H�u�>�� ��l�Wj�B�'z��F�J��׀�Ґ�So"Tvg`d��-e'�!�(�/!��Pg�u?2�$}\���7Y�򓦶N��`j���{�O>l��z�E���b��2�-0X]�!b�׊D�E�e:t`@]R��/�\��o��X]?���;�c�2:�0�b��ˡ�ݚ4���k
	��_���@�+�� �`�'��8y&jB!�wO]p�(���L��_��J�J��X.kf�`�� �p����P�ud�r3��e,�,��|*Ў�53���b�4^FdH��x�3���?��'���]�"�ugf��w �M,��4�C��,��2���q�Ե7�E
���;�dA��R��:�����Դ�4��X)������o̶PK��Yl��p��E�=^��呂ē�H�/�V�#}�EK~B-�-D��l*��B���4\�_c�	��Zʙ4%�!X��G*2j��t���i��_�~SqS{t��0������[��6=^��D����R����$h��k곌m嶖�ksCSٙ��X��
�@�.st����*�6=B2}��	,
��S��S0=@iJ� D��Ʈ��� ��F�Ϫ7�_�V�/���L�#|���wJD:	E��ȑHʹ.(�h{#�yJ��Vii�2c<���� b���u�愈ڗ��Cm�s�t����S���*��(��ӵ.�Ts�&��$���}��Kڋ���@V�z2iPxCx�\�4�t+%Jd�t���۟��O��,��oMS�M��K���.��G����=<�~��Y�'��Ws��QU����5�Uᗶ���2<%:�C���7�PAKdQ��Y�ʰ�oA�w;j:rs�Ä�51B�m�6������d}���E��Y!�Ht�Ȝ|�8*c���c�B�B�Y������b�w���b�%%�������{����Bq��R�|��=1�}HmR�Jv�)�� ���e��\	|�_�^�I��BsJӞ��[j�O*bl�K^�	�0��a�P�Le�1�I/��sI�����^�۶=NL�x�ሾE'���?:�D��CE�ζ�P�fK��]�ɖ��{HGt�\}�x�PPWm�q��9b���䂑i���`��"ࢊ�d��/m%]w֮�H&��<��oS���iʩ
l�Y�2ly ;;l�=���I�f�u"�?�O_��,J��0�i�t��M{I�?oL�^�u�R���._�J�/G"U�I�W�L�G��z^��d������[+�d�~��Ѣ<���rX�O��f�ϭ�7ac��ϝ1፷�q�ٿ��'h�g���[LZ�a�7���ڳv�\��=H��n���@.����N�4V:�b��$�x�H� ��1��c��:�$xG��趱#����+ ލ�T�#+a�h{���镚�X���i!�� >���t��{P?�9Bp�������p)�H��N��z5��W�P2�RC]�랅r?�a�Mʨw���AԒLb�$:�5\�;�:1<+q���U#N�b��񍑣��U���@�+��2J��s����	���\��L:���@΄�����^�!!�Ұ���F~$�G�^��6�;Y=���7&���[�,�ʅ%-jp΍��b(q����=D�,�l�]�6� �g����Y��\�K�	����e�R�q�ڙ�j�o�/PtiEMt4�V�|�2+�G��*s��v�<�K��}���Z�� ��h��:��0)�c��]�R�����A�YQ2��,���觴�C1���r��I�3=��8�Zn��)L&��s�1���S����Qf���2;LG�5����iPC|�5��93�
�SuD�hDg��G�������#)y\jgs�IdrxTAk3����됐�~H��[�?�Z�	��?��錑C�B������`j� ه%�b�MA��7��s�>(@�؊&��uQ�'Ȥ�C3����N�5�S�t;b7x�m$�%�u	���@�ƈn�Y��9Q���'���ꯕխ�u��31���'�&}�=��9^�4����	�j�r3���&��d郴�2<�k�	�D$�>���A]�:�©��������ԯ��s�@Z�q��^{S�S���g/dk
��Ŋ��|ኆ^���}�h���@ޖψ��"�[� f6���z^ިAg����-�X��<�u��ž�;�� �]��\6��R1�!GzO��ff�&�ޏ��cz����%��ɒ���-$���ay\;$3lbY��u������H��x-����ߝ��^/�,�܈3���*̂˿y|��pVWuM�(tBi�
$�,&E�$Wվ�ǪNE��0?���8Mv	�����n��}���z�"�*��.��9��U�6�bzvWy7��Z+��Filf�f�U۴|X�2�@�,g�YR2�"ng���3w�1��A��{��AC�D1a�s�ը�a��d����w�n��ۆ�Y(|�G��r�͠4��@��;Hɵ�E�odlw�>��:(��<��v v��K�r�s��Cj^��g��[e]���Kۙ�b��������Q�������i�)��
�+�Q�^�S9��&>�TE��AyҀI$���$x��%̜n��$���2#s��"�Q���M�)ҩq��`�/y�G�nj�1������r�E`�`������)w����r(ԹZ�uhB��x;�~�mQ̡e��Y���'�1xrC!�:s1:	��]�i��CT���1f�BG�uB%z:Y�}r}��ߦ�8D��Vtt5WM�sԠqx�W�n�9�SSm���%Y!��Tv��}u)3	4�N�PhX��R���=H*�
���e�N�<U��^!��4�<r��K��װ�ut&r�=�g6sY��}�۶%b��]s6+]��)��B����)b�����/[�R"�`�khH;���=e�Qݶ{,�AB���z�ON���͝���/��gP��I;��#��g�U/3c}n@Jd/]���頙,�b�
�*�=�i´�yYϨ$E\8���L�i�����¹�]0\��/k޷��N��	�)��l�	��X���Fy�)8Wˮ���(�C�\�_����ω6�������O��c\�z����*]AO��s��%�j�'QsQ9D(����U͑'�+�s���^���|����d�p�,3O	;�cl<t!'��_ø���=ѣW@Ώ�=�'޿xTQ���p܃U$���ڭ���c�cE^|`����0�TJ��P�~��ʕ�0&�.��~�9�e���"L��u(�t*1Gw<5���9�
,��1�������V�G�g�FK��!�QA�s��L�=U� � PR������=QU�LԤ���K�E�p�2��~�S���}g������qP@4�~r�r��a�:�/I����4�.��F9ޣ�0[<9=[����lbCX=�>�#,�����C�/jKi5L��3���ʩ�M@��`�"��ޅ�"|��ҝk��HO����1�:�7�;�p�Ό�@���jr���_Q�Z9}yZ�:�߁�k�W�,�(���56{�O}�����j4F��H0�n+ܙ�(��9ŏ�:��3	�⏑���4oC����E�Zj
C�ޯyK�؆k�ad�-�0.�^���=����)�:-M���-�a�ȣ~�嚼U�)��x_���/�w(^F�'V�C�qEG���"�����u])���k�5<j�ͧ8��Jߤ�Bš�BA$ǝ�ǚ䣬���x<�Jg��0w��T��^^q�}V9�!�`��+|�\�	�imD-Nır�$�b��h�;ub2&��aDH�(!a��6�?�:���d�5�
��t��p����_�h���mw��Txz���@n/�=�e�zR��;��_��h��M���γ"�S�$�I�%i� 6?���,wgrEY&�4���>Ηo�����I5��6@mQcW����3S~a�Z�\W��t-8�����ύh8�}��<[H6���S�߱����&avY��=n0'پ�]u<el�H��E�PNe�v��'��:]#�d�d�|���W��T�-p ��~�&x�w$J����.-���!u���S(�A���H��{86�֥�<���D�"�Oͤݸ�L5g��������׍����ԉBN�[f��Ի��8>|�D]����.6`0��cˋ��ۓ�pH�N���r'���/����znb61s��j���<���[R?�%����]Α��:3;y�P�yr��R���馌!�?���W�(�Z��hn�
ˍ��!�9�W���s�GlcP@������_P�m���0%�\�K�?Q:,��+f��9�g|��i��9��Qh�'������7�n�9���1�j�CPj/��& �T/�r�a;�j�N��C�R�+x��}��ހ�ve�QN��8�C��Z�D���s��F�3F'$e�T�H7M��Cʈo��z`�r�8r���B��.��Qm3�g+p!�o�^����b;d݂<�4>�CÀ��(Z}[Nq�}�b�_f�e�Q�K]H`R�]BO��G��箴�'�YSsG�d�לs!,q�N���V4�{>I���x�_@}R/�9�xCDUX����D�i@�KV�b��ə����������\~G������ԫ��bg�:��o��D����	�? 1��@�ۋ�~׍�$�i�;�(�ܫs����~��B�ݵ�Y����@���!�S6���P�	����	�E/�2%��q����hy�p�7����e�b.~���TB���yV@���:?`���Q��.$8Y��~��S�Q�y�7j�l_֕��]���c�,0��e@SUkAo$���q�#/�c�3�O���������
�,|r�z�"�%����k�]��@80���_('�����	F
����	h�	br_8�Z`�X��wBY��j�;P�s�4�%m���~���	?w����O��EǄ�1"B�6��h��pB�!8�}�ۿ,�_���ۇO�� 2y�bS�C@V�p�h���OU�&��Ea�f�3���m�O�����Le^I(�Տ�j��T���.��Q����NT`�%bÙ���fz4��Rvp1yt����`l�ޱ;'�i�R��;Jƽ�?�Ы�����i���E�%��M�J&/�Uup(QzCv�U�-�����İ�*u}كfwx
x�(T�_(��3�r'X̤�g��|�kb��[���uG�����mP�Sїc*D@�R�m�UY���� Ӟ�9dU�򶒧�0�*y;�d�JА�9o�\o9��V2!�z��{�|�#�<�^N�V{���x�Ŗu�s�qSI���S3VR�
��O/l���,g���TЍ�UϥWT��a�G���5{�ڪu���~`��qs�0�s�9*'>��I�&�`9>��J:�'E���.$��o�]�C�na��T�FR� !�u��r�Q��B��.�aU��n�*���ӿ5�5�U�(���	L�v�&��M����g'ic^y�	%^���6�:�Z¿N-%UBp/�|�$��a��<q�m�W���:����8�sޒ;?������J�7�-C�+B>��0^�є��P W^s�MĕH�����>!�y�\�.���S��bV�����{d���QÕ=<���֕���<�Х��ɼ�G����nɳ��O&(�q��AJ��
���42��6Z�Z4�����B<+���~���a@Y!����-L��\�͇����ə�ZJ�\0,x[ח��nݡ"���g<�[��1���+�0*8Ǌ�Δ���e�Db�i�ȿ���ՑN�t��E���w��$~��Q�b1+8{���k��=�X~W���=������[���P��A�g�KB�mMr��n���
�����R�j���''�8O#����)A���.�"�9*��~'j+�-��L��аFg(�j$���j	��5�Py�ʐ�&=��~�7��#��y_�El�ዒm7���)�����P�^|�6�w'p��8`B���X.��)��nIl�	�d ^hP�~_³�5 ��5d�E��`M���z]�V�h��;�ި!��)��44���d�Mx�<��:�,���;���_��1ĮTpN�(?�T�h6��
�IQ?��1۠o�&7v���@Y-�R!iL�V%m��`е��#�:��b�*��d��R
"ӌ��=-\���u�������\���@�IL��;~���B���� C�\"�A���v@�j�e��3S�nx$X���~D�8� 99祿�"�"��L�P�|]<mR@q�M�]M+��N���N���ɹ���i'�-�+��YZVn�L�V��<s�N[s��n���
Y.~�U�,j*D��i7\��*��>�(w�Mh��K(M�����i��H�)?�c���C�݆�\ ������]��������Fj�h��&۟7 !�ņes�'	%� ����)�Xy�a�|�(�5��b�2�q=vA��|���e��Oӧ|����[������*��9�hjf�b7�>ݨS�{�4�2��j�����#´�>�5Ə����@�Sg`����v	����P>�
��b�5h,6������Nrb���4?я~qN�*�����<��y��������Y�� ��>Q�e�f����t��afZ
�=���� ��Ev�e���tqIL�'��3]_����8��;�mj�豮!3/���*Q�KS�
�I8��S�!`�?+���C��4���1�bB7R�(PC O����4ӿc��9��Zx�����^s9�o��e���Bܤ↍��H�Ɣ���L�Ō�K%���K\B�gXo��a9w7m<�R ~���0Q��\ޡ�!K�s W����w_���yL�q��G?�2�J9o�͠Y����6�����	WE�_��s��3l��Ņ�jIV}��e��O��7λI*h~+�^�e�� ]���t��WU�~z_f���)7���	(ٶ)�Mi��!)����+�.r�װ��*�.Б�>#�,��1�$N����C)!B�B�0Y���J����'b����g�z9_���V� U@�.a�i]��xiZƕX9#�&Q`(+8���莔��qv�߬!��7�K�ʧ�2Ky�\��1v,8v�$+���'W?&�z�5��QC�,�;&����îyf�i�Ձ8|�_N�����ѡ������^I:�MP�NNX� ����a S��H���"��\gU%jۅ-�\#c����憵� F�`ؚ����\�t�x[M�~[s^�5)��z\&�GΔ!�q����S���Z5� �m�1a�o|�� �ߐ@�t�ALq�#��>rpDi�Nv����2��9D�6d��8N�o��'q���i'I獘��rG`���EN-�-if巵��O�*8ky?�bjܪw�<+7�0���H���� ف`V���
ۣ%jסKe	"�:����~��5V�-z
Һ��]�Iѱ��h*Н�)�y��ߡ�O>�e�5�#bĸ��R�jB��%F�M�]�+�IH��`Ԡ@�Qp���hO��wz)��x	�Uu� ������&��`S�1A�l.�k.�䶖��h�b�qV/�H�V"�l����
�ݹŢ�v� I��.To�����I|�1�Y�J�\B+F�HR��/��� Cn]Zs.1/nT�P��(j�B�D�B1�^��+�v`�`�V{5�}�	moKK[J'Y�f÷;�HZ����-�mՔ8^wJ?6���폂��:�R�7�8]�Q����?̍��F���?H'�/�ZޘxAF]�u9�H��;�=�{����(�l���!�Xi�t�����M]
�M6R+�_o�܌?�0E���r��h	m_/H�7�a�;`�B�*�ZII���K���ep~Jz�.��T�b%�W)�������a/�R�f������Q�Ч���Q{����Q�c�>/����.�m�Ѽ�Kup��������r�0\�Ύ������_+�As��~�݌A;�TB��p��~�ZP��0��%�P����v6�Sۮ���n��&%�{�v�s�hB�ϷHO�i<>.!����@�J�*�	OlJh���W>#S�,q` �� z!��Ԭ��:lG�6�[y��>��SP�}0��Y9�@���/#��:-�`�k+v\X�3��^ǈ����#��.���`�:�x�Ѱ��\b筮�+�9m&@u����ޘ��NO���V٫��A��QhKof�K�QoJ���PKl	��QkU�Ď�g�:�2���,u�U�{�V�͎d�ѧ�`��\J'E�U��.��$j�Ge�����Z���k��0��4��.F�@֦�afm�'�c��E������Ƣ�y���ȕ���ԘYG�\��іM�4�Ø�p˺!������Ɲ��~S�\�zU��K��W��/J��#v����.�^/�Wn#I
oX�D})J�>�+��4�K^Rq�uA��3����`�
4k�ٕ|�Ӯ���Ո+�ZV�2�9�*���,��E8E�����|N�\��DC>�˭������"�#��Ǡ뫢v������X��#�K��Xu�Bo�N�>�_��]�u��������[S��7��z��ң"0s�?�4N�N$0o �sW	�^�w�6��c�r'���S7:�Qz"q:d���3����Օ���~�}��`H��:+��Dfe�)Bv�i$%��.4�|�i��+������dMѡ�ߒ�p���.����t�6x�A1�����{Clrs2���ؐW�U��\:ӛ��gۢ���=�QOX5�
9g�7�DxF��]��qe���v���E��tmTT��is2�W�������AoS%I��E�}���LNnRK:�s��r�@[�}+d�A�B�J(����qF]2?[8�;%���[?3��z����*v���Sq�J \x�ПSu��
	�K���oN���,��Δw)� �c��0�9 XR���R�N�5
����ȏ��2d�ޢ���y���O"����c�G�70`��S�d��m}�U��W\�����b��ȉW����r9�T�I�j�I��K�g8{#�  ���rI���1�KT�K�,ywHT>�{���˟LgZ?)��W[ r=��I����)��,�;�P�y���U�gY��1)�ܞ��h<�U�g��n�Twei�/���D��W[#G��^#�dAE~�3u���N%�1\�z�y`Y���K�nY2{w��Z��%�� �mMV�U���!M��\,��,�˕{r4��KJ����k�h'�݁����uܰ����� �$A~ȊpY���$�F�0c	_B<J�td��J���_����9U�er�zO�d������N(�r�s{cM3�]��Gƚ�ƌ�7�W��@�IB��/�$y��M��e� ^�V���ڈ��-̄�*,_y*�����Mqu�4�|z��^�MJ���XOB q8��\�H�Cb�uˬ:Ƴ�JQ�JT�s3���V�S���̶��^ǳU�������5t>�4��z��Je�����H���L�İ����$�iB���,���^ۧ_��N����
r�κ�v�S�f�7%$���gq@�������I��<�x���
M2=���=j�� z���'�b�O�(u�v<f��(�ف�4�Ds*88N���٦��^��=�a����S={uw���%�H�3��SѲ"�uCX콤WDF0�85q�?�Ԕ%�h5�ɶMOr���(y�8�8.}�1�Ғ��>g�؀`��!�l�%-ǹ�,�ɔ���Qr���^=�9Il��J¡���V��S���
��b���C+ؠ�	o�(�I,,��8�ٽ�5�������)�n�"'J*S���$nM�еk�����dE�L�te���q�Wx�Ӕ
j���$�$}�LO�æ��;�NDˊ�ұ���7'��_A�BV��3�<H��Xr������Wh��jQ�u3�9�v�(R���^W��p��.��]r:��,��e<뎀V���&E��9�	���%�����|5Eq�dv�	ب��p4FetϹ��k�,^u��`���ju �y�$P~��\�Q��Օ��;m�<7�6����e��7��0��l*O��#e_$�w�b�"�k���;�w�o�F���ɳJyīE�b�)h�W��8P��vi�Yޔ}h�"�6�����l5A�\Ƚr`� ��k$pj���Mj���f{�4ԴQs�u�R���Ɣ� }c��@>��S?�������=���H�u���+[~�%�G��N��1�n��DT�M|V`%��2%���Y%񟝹��@WJ�p(np�(N�@x_��v� ��/�����7@��t �W�������W����w�㨿p����3ێY7P��� 9"��f���v�@b7<~H>]�Xa9����9vq�ͭ��hY��^�1����E��nr5�F|R[��,�3͵�IHN7�&���{��ό�C��pղLf��"f���x ���~gwHo<�´�g@,�_��������c�X@�_;��t{�9dj��>XT f�����
󯀍5�ݤ2k �����!sd��>���r�++��$¾����g
$1BJ^]-mGR������d�B�z�ay`b�D�Q�L�@n+�X�y��x�>V�.B���üH�l7�pb���7�@t������7ZV�̠XPo8��Dr�Ʊ�J�,^:d��$~���?5si�ᶻ�S��Hj�\�L�A@/;����+��ax��Ϭyi�/{|&~vNl��$�|���Hk�@���p�b���b���3>y�� �.�a��.�CIR�3ԙ��J�|j^���m0Q|Ť�Δ'��sN�W�m������q���ɿ�=�ͪ@�sg��g�D�߻���B����r�'�z�>x3pG���r�#�W�vOϐ�	��c{ƲX�4ƨb],��q�ZC���,NI5�C��Ʈ�o��������u����������ol��o=��2��H���KK��6�ƍ��1�R�'v����ַ���f�`���m��y�z,	���^���mW��[W��r�.�+��s�W%$s)�����Lk�����°�c;������앤��8b�VY[��v�����`;���A5,f��C����~\�b{�`z��с9$����y�qV"(��{�z��14�&W�S� H~�^�,kRa)k�'6��\CL��WÖ�
�J�������ei�T�"N�o>5F���#���1ڈޒ�n��,�N�:*�B����Z���CJ�垅YY�����y�`ٸZ�}�浜_�-���2���>Y}�LS��&mZwF�x�8R�|-�_�Z+���X]��f���O	�8��,�T���(a����^g�}V ���|��TԎU�#4�����a�it�N��9�����a��{�F�K@0Hʿ���m��|L�(��U�5�8��t���靴��kX��v���2�~9�)w'��8럾$*��Y��mz煮_V0M��g~��5�ɤ�e�O+�p��"eD/R��%�O�b�ʁ'E��UQ_S~{��=��-$�������*X��gBe|��h�F4-��Lk&��	�>�R��{೾B�g�H3�X�?�[4��h�DV���w��.ɮM�V_ �� 9D�j!�^G�%�؅S��u�4/ʚ����^��p����8�Sk{��S[FJ�fG���D�1D�L����x�]ᏴK��?�'4��N����Y���;?eA�ƴ����܍�S�1
�5K����A}��E3�e�!������������5sb㔭�vW���Nt'�r"n]�R�!��y�,���
U�b��Ool`�{�8b��F�������e�f�P��RN�@qm��7�¯��rY$ � !�¹��S#�����]:$����I�c�6��Z�����s�� ]�~�(����LO��mA��=G���]�Ȩ��iJ$�6xve�M����ЎE,�K+^��$˗z~:M�h)��h�������ō3<�D��L��d��g�2�]~��Q�	9��t|���H�b����,��[ c�1=�?$���/�q��__��"袷���bAT��P}�)7��[��U�:��߯��n��n�v��5|����ȷ�1���Y%0C/Ĭ�bB�=,����'g�������G��c-�c����/��I��r]�G�&Z�h'��m�.�q�N	�M��ǛU����C��1���F�aBJ�Պ�������Y���ސh�X��p�q$|g�/F�7��������=?an7����?\�I��s�����$k����@���v��b�J5�dO�
T�QQ�F��YpU����Ijad1 ~��,������}͖|�
jX9+,��z���\�+Kd�pE����̊���U �Σ�����g/L��Uңہ�z��\�,��ǧh���� ��� Qlk�|���
l�
�����.z��Bg�5���?�7����bPq�8xU���f�_��
���݋�ƀ:����+�HK��a��lC��_�JY��~ě�ycз\[�C��uA6������ß�w-���F���8���h�-kܬ��$Cw�[n�#D��M a�Zm�E�J�~ՙ��=V�b2o�A1��L�(p�@(����De$�N`�������m	X�!8�m*J޲IMNE>�5�D�B��M��x��x�'���&&��Ol2�D��ϑF�v|JT%�t.��.��+�]C�|�S'4�:� ����`�C2~Ե1���D���[��0ʛi��[ޘ>����p-��s�M�`b~{������k���0��}���T����ʍ�S��m?��[�X���C�#����UQ
��xk��&�ι1`X�B|M ���d.��6%-խT>Q/�L���|��?񡮞���n����΃%ŗ*�ʿ�Q�.�Hp�pm����C�Y���4�S4�.��ƽ���F�CkH1�[qI��2��Ϯ�Z�*r�F��Z�P��W��w�%�JGl�.�c��$1�RtQeCs�v���imhk�����$����Ԙ�H��~x�*0��PN5�[�ݕM5u8���w��y;'�~9�o�h��[�8�����t�5NES�1@���F����`���ܣ�o;� 2���\;��.��tJ�P��g�㷭cن�v�>�O��OK(9��#s`T?�;}`�3����殮����Rt���3y%��S��hE��5ά�+	^����л`G�.(#.i�C�M� �b��� �QPO�{����E���� �H�\vǯ>�Ya�~�\**��&�Th�����>]���a�a��\�L9ˌ�&��7#�Fe��J����A����+ط��LrMA�t�u;��m<¢�U�/W��o>+��H���6�������;g��_�F�0���>�,���6?Ǻ3^�Kʋ�� 0CŶ�$䕾ZQ�K�&��(�FE�L�Ƶ`ߠTH��N/8�Rͦ_s �Ra��5���L���g�L�Dl��6,Q�Y���P s+PT�oOq��"4'�K%�ɳ6�)S��Vծ���uf�r�' �_#=,�������"�������b1v*.-�o�]t��8�a�mb��Ը��=�����_/��TR��s���20}릣0d��X1�r �4�>�� �|ɊD�s4#5x6���Ųr��k��(P@�����q�5 �pM%f�rt��I��
���I�>��3W�C�ںe����	/^%u!��/}A2�����>��;�����wn�p�+w6aUu��m�(m��A6T�����3��R?�PQ�r.���<��/�C��bڭG��Dq�*2�H`��w�
#q�:���hR0:��T�54ڠt����,DQ��y[�:��[��{�^s����?%��Np���
cSz��i�~�V'O��$8 �J����;�-�J�����.��F���U_?)b�gV�sZQ�P���=��^�h�P�Q�Wո�<9�=�G1f&ų�-�o �2��#�_��ң�k:j���u��,�'b����M�>�&Π"zi28O�����>�nŋ��p���ƕ�� ߛr=:ߛ^�CT����id�6iE�+�P*�pT��6�$�Xw��ƚ]��+!�x&�i�[ ����V7�;�Z�j��/{�[p�W��zY�ՠxPmC΋�dF@�h��բ
O�؇�n��|��xg F58�L�y�w�8��I��6��h*�-��\Y  2bQ4��tn�o��66�<i!�<T�\g�����U7VEb�zi�
s��J�jFK�u ��L� q2)�Ɠ�o2�耣�x��n�3��T�۔�6����'�������5�u5��b�tD���J��L�~G_"P݅�����a(;$��*}��R��� -�ij�5��B�ӯ��!�W��j�ہ{x���3��V�Y*1�2��O��N@�J�?���N*Kz�e���L�~\���a��&6l0����C��+��>�[&��X�7��Ӗ�ʙ��p�<�����gu.�_r�ް���4����d�B�(���TI�,�w�2"�2��تV���ƅ�6�2��aq����L�F�&���xRd�S�օ��R���I9��5T,��\D�[��ݒF�D����Ci��2��Ǭ�;{�⸃_��ÿ+���.��X�az��=�;���]݁����S���J:YkDC��2���}f<��tD�t��l?t�Z��M�~,88����p?&�������!1����>�!E��@N5�I�u��i�X��1�����
Ycr��1�1>��������;ip�����D]�͌ƺ��n&|�t�#fR�W-���a��(k�W���B��@�؜r��t�ƾ@�ԩTE����/�G-Z���� ƜG@AE�����a'�w*#^�2��|Lڔ��Ъ�T@���1�����ot�T'��0���樕ವ[� T�#��vK�4�e2�a/S������!�t��'i�[��Kr��kq�*�l�r����(OMK�\�H�<�r	!�*�
��?eR�l���j�8n�>��O�����}t������hI)o$Ũ-s7n����8gݑ�0'��q$��ƞ�x��ۥ�Ao�[���Nzmd
�ߋ|���u���`�8�E]���Ә��7���?�� L]�����T��gv��7��{�:�pD}�0;M��	._e@�^�g�lI�!�'�8�Zب�DF���Gh4F���5�T�֖�Y�?��>�j��Cʃc
x��|ћ���d�34[���aG�{$�u�\cd��%5d���E{�~;WC���L����Y�m9R��T���.;E��RGL/��"�be�"-��P ��,�:�2b�ߣ:�v%,ڻ��_��vB����Q�4��Ȥ�t��8����Fg5t~�~,���"=yq�z�����d���n����<~� xR`D�iy���Fܡ�iA)M�F��@b��A,b����ΆkQF]1h�K�d��Λ��b�.}�+���+�A)!��Dm�^ŕo�Pf.��4`�X�0H�D����h6#� Č�^�tp�l�k���
S�_GH���sm�t�Ik���.�TU��\�T�j�F�$��=*�������
����%'e��-Ɇ �|���#a��B�i���(m.at�� �[����J��dF�el'|dc������`c|�Ӷ�3���-~z�$��21	F�,��ȳjM��1����Ɠv��:�Y��[�G�"7
���]x���n�ъ�[�G�S)WWv��eΡr�7�8[!�v�Ͻ '�����pP�B�-��2KP�}2yR^�y�2x&��4�g� '��rQ���Htl������q��ǃfШei��J7v��!�w�С��!
� 7yH���ڡi���d�SKb�`%��4&Ҟ��������q�Yw�T/����ř��Wy�`�Tϕog��^P�;���L��7���Y3�yP+W�!r>�J���7��`ԡ�a�E�AY>��=r�Ƴ��	�Qƚ��(C�D�t�w����V�#����I�˨p>���Rݲ4�~��C�d��� %���%m$O�ig����3=�m~�4_��9KA�����^�/�����y�����	c6|��*TG������Δ �����"��{2������XaS�B�_J�KS%�(��A�j���^Y 8U];9�@�ʜ涒3XX�M{�޴%-č[���+tZ��G���ר��$ߦ�H������Ez6�rP��oo�2q>C�&*;��]Y�ɎʿO�!�3�����H��Rҗ3%��`��:��L�H��J,�?�ڊ���LK~��=D��uC��y􎓹� D5&��PO������;G�.�ָ�����վ�f�a�8t��?�z�������m�ǚk�����I$���$�J�ﮰ��#w���s��ʁPW��R5�s�is֗h�Q��52�G��{`+@�¸:��
�9n�q����h�tn�;j�X��%�5�U}k��F����g;60�E�0v�J?�[y�������V�7zE��?6�fr8Z�Y� 1f?��ϣ��5,�S�I�'b�%#�^g�[a�����A�*q� 5�j:����i��Q*�w�$qH� ���Q&������_�\�l�7��c�J�<������?{�����c��Q"
�ňTՃ��$p4���;�h�-��9g�d.\���F|";�(aM"q���*Uof<Ԥǭ~8M�t�1��ߐ��|����e����<n����n���ݖ>�$Y6Ԉ)�P�ڊ��t����IC�R���ML$��gs@��D�g�+���,��^�����˷o�Z��釱���$`�����\���$�{�������:43�^<g�8��]�xg�5���:���n��u���ro��CEp	�*m!/�>��Ѫ����Dq�Ts?b'r�����{E��,�����'����ji����`vِw&.�!bBBu���ާ���G�CE���w %[1^�nn?���ۉ-��Y۴4¸����58'�d��������+�A ���&�76L"[���*�?�v�'z[�5^��)���t�@3F���1B�*dV�^�P]̇�'wd���}�Y2B�M�y)A�|gͥwn��;a"���
_.�4���}8����
�.u�Ա�m�v��D�b)���;�]�h�ͬ����%��M�֮����='U尀����j�� �Z�q/����tߜ�2y���3�&�j������و��q�����&;���N?R���V��}׃Kݞ���}I�^��윤�E�R�sz�|���X���l=����2�:i��cc1I�N>�D8�;�,4S8��$mz��qsu���ߡ]�g�nD�<SI�fM�.�iImϭ=�6
*�!L��v�~�5�2����i�_S��)�SE^{� @K�m��y���+vne�m��=5���4y2�T�}��XC�n?�m�9S����ON��T��(�?Sr~�*e�ְӸu��|�Ԡ$SX&8�j�����P��7�<-��ؠP�,�X*n͜k�֯��\C�Ͱ�i�D���V����|J������-�J���ӯ�nY��(T���t�Efkp�v��R���������k=O�\C ݪ� �/�-�p�
� ��S�)Q��E�\k����7�noXl�
`�>ZO�3�������A�x ��#�D75�`��D�l\;a�PY����i��I�z[��e�fx�ȃɜ�xy*c$�aSvE|<t&PG��m'�� �F�˻�\=�M�ƞ�_2���*�5c�"s#�f%�����VЩ���eӗe��:���^�s� ����<��?�,4�^u���:?D�k�J_@|�Y1<��k��ν_S��te����ɩY�<�-���eML̐���	�B�3ux*���
ɯ{	����G��#VC=��J��,�*6���X���:�����YCP��׫w��n�j P�1ɫ�7@�4T�fB��H�/��T���]P�!D2a�S;E�m��_�#lp�&�,��ߐ�Jd�hQ4�p�S��+�eւo��`Ԛ�	F�Rm�Q%�}*�) ��r����0��
�}�z�U{��x��D��9�#�!��P�����>)q�7��!��-YR,���;�u�8�6.j��C�>��=r���U��<4��XME����qތ�;V�Bj���b�'�yv(�*��n@UY��EGg?�&JO��f��o�id/_ ��(�2�m��Qy3��B��җ5��� ��F���+)W����G#�s����d��E��M�Q�fG���������3Q�J��Ů���3�y)}���X��Sj�Րs󙉹��g��+�A����Mn�m�\�@��D�{�V4��6�"U W�5K��g��5�0f=d��W�l`��D ��~ɀ�G|�,��w�r�+�>�[���p�VD��L�bi�<E4��N�+fJ���!�U��M8=�4!D�^U�U��?�z��'���]4�g'�#�8��8��_����%�J���8]�������z�I!�d=���dr+�$�������|Zo��5�B1iAA�뇯f�7�k�	��!>sn�!o3UL��5b#��DD���B܄I��w�L>��o��3q��y��P�8�����Z*Vu7�d�%d�ص�����-0q}>����[�l����&2�J|;u��}Ãf���?�����(x��$��P;"�1����5�ҼcLxK����fZj��v�9e3r
۴�{�򭂇"���"K�@�@�1�{�5՗pa�Zn�>se��Սѡ.v�j����� �|J�M*��v��fu)i��.J�?٘raߪ�8��M?�=n���ˠٮ@�)�D��od�v�mO�q�űj��+>�6�Д�
��Yj��4PY�D~�jNGh�,�:���������N�f����ƿ|ܔ�>���j}u�{i���)�oC���sQu�E�o0�V�#�����;ʷ��:� {�{:�hB�	Ѽ�t3]����U��A_@�������@%)e-O��h;3�� ����v��#�X�|Ӫw��ꇎ���X�m:	V���~���Qq����I2��w�n�I��(E�0(ٖ��� ��{�f@�,6QP]���\d��g�c�Q���j�՘[�^
W�`�P�d{�J��0YR��%�\,��"�BN��5{[���U�H���}�뇙$(����@l���5�EѓҮ1W�Sם���a+d �%^D�#]i�@>#UבS6�����%:�����A���� Ƹ Ѹ�D��n�^y�����FS����&Ĵ�����ʐ"�A$�%�$���5��H���^�7���+B���L�i���j��\ugyd=���G�iܵ] u.4������	6�v��O��urX�&�j�P�:�~��p��i�'b��8�g�wkK��3�<R�;zw4�y�9|skD>u'�-5���%\:�(��R �< �"73��}|�KJ
I�+���G��Tw�K8ăsJܲ��-�t�o%n��S1��)wI��^E����MZ5*���+����]EA�j�5�;��;-�*7� vBo�l\V>���Q�(���Xe�\��h����k<��v x(�(r��N��v�}
����5�]���imGT���Ϥ�?3ϐ�����'V��$E�ҷ�_e�Q�k�i���A��;,��y�F=�{�i]�X�־ġ�1��0o"߸~��SF���X�F'ΟV&��R�P}�I��,�Z���ҍ��0B4z_qV@����X\��:w�O"N$&ך�mU�0y*��=�!���W�i�g���xe�lz��-(V��lm-M���qZ1n�v����01?�z�ʻi"����Y���#<2���齇m��w������4iT�|��S(_�q�W�����q��fn��zN<g���`�.�w��X�q��T�K �\\�]�>����`vHv�^��ۊ��?��M؟�zH~��7�{���hq �0��:�}>�M�ik}��F�* +u��)��ˑ�p�~��L�����˿Y�'("����D�p�X���i�aNY]ƿb̽c��Da"�.f�V�W sF���0��1�����5�@�{e��_ңI�ِ��PV��)�Z@g͓����VP�tc�ڰ���L�Z9�r7���m�ȚC'�e���?��7�7��tC$ĸ�� 4� d�-������%��;M�^���i�-pW������^�Z��_�jjw>2G�o/�D�����A�n�j�P��!'��y"aUt�w��?l#f�`JwUo��� �S��4>Dv�2L�(63��f�LC�VoL�w����&=�d;��ldNUL|�?�닎�)<{�a� �C����Su�ȩ_�WP���%�AK<CD��n�2W@�Y���!y�`��>��^`�ŀt��t�֛g��#���>S�bq\��"�U��UȀ `�w��'ju/��0u���Ī9���|�s��=��W4�P��,����#1�ۨ<���8&pjqx�ZҒ_�%�|+0T���T�]���;p�� �F�����T��8��[+gU���ô�w&�2G�~��˜��w�K<��G��A�����L�3�,�l��@/aҍ7��M�4q&��\dLh���v�C����Ä��Ϳ6�]=(��ě8h���QI�C���5�F&�r�c�������hg·/�\�v��e���_U�� �A�!M���.d�[y[\����H����6���>�~6���M����F%B{�S-�x����ɣ�vm���g-w@�p1��bl�['��%5C$�x�(��"�wQ.{&>��$$	*�N�(?�J*��<���6�����p��=��]Kh[2ܩ�����ih�`:������X}��M�6��C�(��6�LкTR� �1��ol�2�h���u�x�:�SwdMDjց�#�\�ٴ�q�!-�Q݊�h����AZ>8{d�ezK�3+P<z����XHS/M��>b����e�MK&�Md��x`)=4(�#^�k���PH⨆�F�^=̰g�g�hOR߱W%Z�c0ȍJ`!��� F�
t���S�gL��*��Kױ�&~�k�@��:!�i�'(���K�8��#72~��>n���nN�V�F��J�cRZVQ�K��N�!��ݻ������vS�&N)��V��}��C�?��cf>�>_0u?��0�i��i�ؼT�v��a$�v�6��$ϼ]�7����IɡG�E-Z��j����yY�����0�N��	�eb�I���9}Ƀ�?6�Vz?�yÃ�4i�H��kWH�B�Q��fk(�J�
`Ȩ�
@��Z( �PN��fb�$"�X��)�~�0��/-���8�e���SV�u]#R��ۍS;�"�Ӹ�7^;=rާ80acS	r�8yA͏߬���T^ZՀ%��E/����,uH�(�u�)(���Ƃ���9ȐOW�+�~
�ښ�hbQ�;d!=^��o���*�o*޳w߭]+�ݻ}�y���-��LLy(ּ�l��8�7cI�y,9�5����P�m��
�����ihLG��|�)t3��e�\@D":(!d1KgKm��=N��!�A\�Hx���#�:m�_����7� 7�KD���w��>&&�@_k���񸮓3m�Y�iǜ��XC^���J�%��Vv"xE?��'3� ���<���"�4�=��/�2�������JO����� �UlA!��T���.��|g�|Sx|��V�BR^*�Կ@�&�o���N#w�K�MbYn�Oc3̾�k^����A:�xm���dk�~1�h��r��
��k��/�Q��F�f�Ө^����?~��Y�ȿ ��;�+�L��l���'	��@i�f梓?��Y2cN�4|��I�&��p4�,�B� ��VG�e9W��B'ެb�̚�v�_���ۜ�.Gb��:�A�r}Û�o�#�����g���Gͩ����Q�q8m��qԫ�Z�U��� z[^�Җ���j�B��}�V���E�{|��H&�tDr��.e�qe��o:�ճ�C�DjшU��y��$��+�/�L���6���t]��~{�I1;K����n|��:� �)S}���S?F �m�A���^C��RP2��@A"ك��HF^�ostL!t�����a
�y+1GL'��AN�p +�}��t�Qg�̇�Əc9,(�pe~]A�����R��[�}�Ա��X(
�qp��xU�,QI���ȩ;��f"LdY?�r�\�������/?{�V���������|,#���?�ɽ��+�AV�qP)�""��O{���֜s(��H�]F7@��,��F
;�ޛ޻�o9��m3���]w��uz����w-��9�m�lAhqu���<����~�R�W�*^Q�&.���A��E��č���Em�ý��Q���*�u8$�s*�0֓�<#E�O�9�8���|S��gX-)4s�w���^>ýL�aR�
��K��DD���P�tr����-�Vf�����Ed~E ��Ժ�_�НT���`d�{0/��W��4�Y�;�](����v���Z�E�^�yh������GVO��VL�ͪ�-�}my�.[=#�����Mu�?�eu��<�HG��IT<Z5��B���n{|�9[��T8�9���Nw �S>T+�.�_�8�4:+6ȅ��%�2�A:��b�5YP�Gu%�{5��o{�� NC�n[0\�[>����0���ܝ9�,P��eO5l¦�2�GL���>��Աh)�N-ەU9�h9�0�_�x`�X�*�e�X[�/��z�ĺ}�Ш�$��#�xm߿Ԟ��K�WuR��<{+�
�&dl}����� ${a~E�[ngkS�9�A��ޫ�7b�������� �\�M��Q�o� �K:�,��+.����j���'�S�/��	P=H!K��>��r��}��界E��"i�}�
u����G���
f��Czu$�"���Ҍ6
��\v�.Q�F_+�y�XqH��0]�����oRxB'T�y���(1�t&��j�-��)��+�B�.g�}(u{�J,h'�-M�x>ק{Kn?�Jω�)o�{�0�,lr�����$>ww�P���27���1���MgO�+��R��Ar�.� R�zi�@������S�����J���:X�)��(��<��,�Q	]=���o���焁�P����t���d2�6B-e����glA�13�\m'Eܜ{~�p�Y��_$����R/�/s�/w�� X4g|GZs����J�]�n+O^���_�\��6j�����:cE=	D��s,q��Y����Ut�T�W^ϒ����ɽ��yE/����G���-$�|%f��n���&T�>���'d@,�I���Z�����Dⱈͨ{�ȻiS%�o�'�m��t���rV�� )��`Qr�1�<O�j������ʖ(��p����<"
V�{f
UZ�
B�v��XHW��F�Q��@MS��!{%kôv��u�	�l��r�FaR�~��ݱp"�hٕ(�{�ؒc���r��Y��0>�j`ej�HL�->��z�~)�f7����cW����T�6�����+���G8j���� V�h�:�ϲ��en���h��?Q�R��Q$h�ա�� ��I�V��Mks�6�F���� �C!��ˌ��OX�������Op�,��D���P*d�,���7��6�R�YE�edC.��a�/[����Z����F�7`6f6��:�V�0F� ]3p� �(w��Zw�^[�����Lƺu]�N����.~\��c����w�Fn�6��6HnP�����2*a������=�~|�/�'���AD�&q���l.b��8�pi��g:�懊��J�I%�e�O��Б2��"��H:�0":y�xT�8���gq�Y��T��
$g�Φι�Z���� 1�Y��6Q�M\�_cWT����p8� �~���?͊֨܌��fN�RI{H��yM���s݃	YE�ީ�ּiW#|�y���=M��:���R�w���
�+���&��Rz���Ӥ�����`����݅xLĈ��ʯw	����F9����-<	t:-�����>���?X�j	5�J"ӷ{��WlK#c;[��e2����v�'x�l����S�r��C0�S��[��s�Mg�֓s��zD�&��p@;�F���NI[�s:atb��B�G�qQ�d������z����r�	�|���矾���c��yx^�q}��2�4���7Z.Am�گ���I�1L�k�rji��	pW�������0-zW���Ղwق�l�LO'g���x6���)=]`�����K'�<�\sǺV��V�J�Ү�hZ±�W��VΕ.�v�*�f��oF�(�$�����!ۨ��)���?X�ԁp�ܯ������#�B����'qq��N��~$J���ޣl�p}�I��b0A�TV(�k��k������q�ŜhA�a>�����DmȐTJ�m9�iͤ�I^lh���$k�L�D`�h�i��x�Ey�6f����Q�<)�ދYk�^V�)����ѿ�`��ట:��;`#l�In��f+H��/Ơ�)U�3�8]�V��р6��S$�,��_����F�H��M��W��.�f�`ĺ�������>;WO=��ܳ��hWո�tU!�v ��Q��۷ ϲ�He�|Xo�=m΍��UD��ū�&n6��.�$��%"�;O';����/XH�����h�r�u����c
�9L��Kb�˙'L��]���5���ʴ��� �%(�	-niiD].����h�`�:t��'	�Ba������ D\�r�9�]5u�t�dL�K��d��x؟{�����D��XV8R}��S�����0;��p���k�`\򍸪\=*M�^y��c���\��}��T�o.4�ʼ
1��|���;�����#�G��$��X�����qw��R�S&������0x�*a%G!�S�Vl��y��X�p��`y�_�Y�hw�?1dp�3���������CJ���<���7<L���sL��\�������4=b�E���[@4,�iF'���i���0���8E��F,�%AQu��j8����]��R�D��&Y�x&�O)�
�#���U�$��u;%�f!'�Gu�.���2���4�#�]�n���1]Q�}�M�%3�zNeh��8�AAɈa�����&�4��$��<`�cS0�F���!�N�Δ{�d����at�HV��An'	B�eA[����GA���K�C�d��S��!�i'��Y�<.�, �V�kic-%�o�>^��#S��2?"�n{#X�28<��:��&!Jm�G(�;;W�u-���9'�نT,oV��4�����O6�^J�go��ٻ�1�<8���9!D���U�Y!M |���{�mR�U�'H!�E���͉U;_栣�W����j���E���x��ڂ��ߞ��&��O����E/��U@�j+M1&�s�f��@@�<�ŚF�"2�5������Y�I�����1�ާ����S\VyI/��KhHP�>h|V���@�@������ٔ��!�x���QG��]WK�f�`�o^� �$�<u����y�mb��i]���X�WUv��z^^EmAq��96.�6굥� ���)|\���JX�t�֬��Z�j��q�.d�����f�$8U@�;������"�`dt����Yܨ_�����(���͂v�$w�WäfJqT]�����\�_�E �!�v'��Y�� �z�>�\:6�ř��#��D��� I�J��hq@t�c��I��*�J��SD�3���+�"���D)���8Q-
xe}pEy���g��jɞ'������Ok�o�X)i�K�0�6i'�>�NPNG*	Zi���r[�=uނ��v���ٛac���+mo�"�(��ؔ�ct��x� :�˨ïy�����U�ҵ N<�-��V)<H�N��7Ƹ=~�R�E���Z|�xL�)H
4��K1��=ep�KH
-�����3�"�B����M�\�̃��}����9�n�Z�ϱ�W�ɓ�ƹs�i<Z�aaD۱�<���Q���ۮg��k}������C\e���G�DZb���<½�i4tH���(�K{rgd�>�~,�L���\Gշb��*!~0��4D����Ə�ʈoB�f�3�?E_�_�(8�v����.����_�G�b��s`H�����*0d��l3�D���X~A���a]mb�����a�.4��YͰ�e��|>1O�i�7O���H.�Ħ��Hz�qE����C%L�CcG��;�a�+VY�G7�)���90�!�E��e�^�]>3���>xg���!A4���p:v� ��RU�>��Z�/{�
	�\����V�^{!�%#,sԐ �4_"F�+��H�O�B`���X�.r��,��p�lb+jK)�2[
*��!-��"�&^ҳ�S\�)�-�e�A�ML8}�.�~dL[��1!�@��
oz��'��������E� \<�{�&�X3���������ާq\�B˼"�=�}E�Q���gr%.�q�_`��ªW<TG����L���o�
	K�8ZU#���z��B��ϟ��
� ���M9�ʑZT�؈��=6(��梬�2�9*F�I������V��q�8,6�{ty�Ǆ�#����"SJ�+3�i��_�|�x�@NhL�"4F���`S��n�����~n�FC8z
�=w�>{���CIaW�P�id/���04'����g0���k�ܮ����p!���s�>p(�FT�"�箃�����ĵ����-��l[�<���������6�/ڛ�&���M	J��Q� K���{p'�p���y�����IUԃ��ec %-z~
��%�z�4���a+�!�kׯ��f��P�'�j��z����9�9H�-�Q�`,ثdpa�r�-N*J���*������h,�ӣ
��	˄��z��ZB�0ա�'<f�uP���m�?z�U(=�Dֱ]�{Cl~H��נq{b�˔�uߌ�9;ݰLUXa?���z��B�I���ʔ4���R�\>�-��Jd�T���8�3�S�
��0*Ԅ//(7�x^��r�-�1�(�Q������A+�5-h?�I�*u�:8��L�сV�4�#Uĉ���p2�4i,�Ի�,��n2��t���A�I� &
��gE������<@�"O4fcWiפY����y�WP�Y����R&����Y��+D�����Қ�����@��9��Ş��\ZQ⽒/a�f}��Q9+R?M����Pd�%��H-��/��?i��ؿ�v�ܖ�Z�~��2���|Wj�x�ɥ܊�dJ��D�e�_f�R������x5ɗt[Iw'���1?�eN�����v�e�N yMrj02�]7��ø�f�f�Ħ+�R�D�c>�Z��)%����g\�a��p�
7��Db�{�I��F&����C=����!	�e� �Nm�}@���c�1��$�~`��?%��7n���&h�> ⪵�E-f�p��q�����,뙓tw҉�ap�_��ob��J�ˍ�y��03��lL���b)"T_�,�����.W����D"�%�P{5#�'B�dk �����$/�Q �N�6i�ў�i�ѕ�N��WjBʿ��{f�������$Db�4�ĺ��*գ�`"�y�$1�����&�i}J�b7��G�+Z�8B���Z�GEy���tn�)tS[��������7��7z�~6�I!�Yic�Qߐ

8<~]�ZU2ۭ���Oو�t����:}�n��7o�W�X��p���G�vo�]J�-7j%w��/�Vy�sAB݃������a�yK�S�Oj����7�g�	�2��Lb���%��+�'[��l�j���ꟃ!��iq�P�`ݲ
i�`�JU�^��ov�3e��V�G�����K�QQY�9JB!q��ң�i�y-��� �r_�8�-m��^�#���se� ƺ�^p�1,��	yuc@Z3����K�a_U	+F�_]Ɯ�qS���j�}��_�0�T�P�4��5��t ꌏ���/�:�[S�9
 ��Z�$�2<�X��M�a���k�N�RH�� �W��� .����j�L�l,\IK�al���U0���I���Do�2sQ��L��;��j�s�a�ţ��wv��}�O�k9d@��ƚX�\�hBb��1:R\E����f��±�o�n�����~;˲��aC�ܴ��U,���04x���h�(��`��|*I��6�U��6�>'�~f�DbH�/��_X�?o��,֧��
g��U�-[1���E�erS��+_٦{-SYk
��.3����#^x�u2T/�3�Ն�2Z���@y��h }P3w���DB��Hi`�+&�3��#J[3.f; [#?Z99?��;!|�㨾�9����2l�^�S�w���ߍF�$I*ʙ�H�Z^+��'�q��QYŖ@^����L�ȡ�!q�#e��L���H�-��<8��~g�c��cRARj��W��Qŉ2v�.� ��h׊㨩e���q���jb��Ъ�hh<�)k�`�Jn�Q�����3k��K�4��_#B���Nc��м�|ĥ�}�!��t�'��l�W��P��3w+%+�W���Mr�E6�G����OH!�������'��!����`�塋QT3:�:�=Iˆ҂]����`#�u�����9a�#i�@���d�TU��k4����O^^���:��@s���X�j+�9٠�쟸�:�@%��í���kI��J(����MU�E33��(vJ��ա][,��4i�7X}�\���&���|����F�ڑ�������ѥoeO����Ҡ;�mMM�����F�l*!d���6�N����o!`��ӑ*�c��Bj�V�;�Pje"�u3��e���T�S>��9	�
�9���ˍ�g�,bc�M{o��#f�n?��y:難��w�l��(�J���)�w���1~���X���~����WӍ�؅�^Z�i`G顴��7[E��E���9��8�����`��~|W�;�p��Y;�l��H�U��>rn�ד�����lD�\�t����J�n�/=��YOE��0<��������5�
3����b?�{����x�L�<V7C' `��D�1�0��龠��b����@r�M�i�]�;.#ǌ���˪���V]��ꊐ[�9i�]�cK�/����������܌G�L.�����8�1ĈPNo6F8'����\Y\}�y�U���m�`R�'0�s[á���5ޞ[�*_��r�X@��,d!2L�R�4!p�~1��`�v�_��c���Dw��h��J{4P���"{%�[���@@g	'q�P~�%&��ZD�؝hF��	�C���ˑ��8��%KBf?c���CG ��Q._��D�z�)�fX�*��u���~0��x�ݪ�pX�0�{�R�W�0��l3��p���O �..B�	��rŵ�L0s�]�`!#�&\c��U�QZ�%���El�
��J��zr�y9dv����D����v>�ڌn���8[����!��C�z?��JP�����3���<��}�D��0`whv��1�bj{��P�n��O�܀o�NXvl��j���3�����&f~���og,�UX��_AWƏ�)��(+f�Vt��Y�D��l�i`r�E3=���C�(@�']a�>%�f�U��o`���m��˸n9���^���������wBI5�%w�=�/���n�u�8�M6�����<�VT+\N��o�ax���$:$���¥�A��b��{�S#\V�k��.���c@�d��
���!C���Dk��U `�?�����J"rVǍ�U\����C#& |�q��)�Z��/u���!D�(̦=K+��+�ڬ�un00�b�H�&e�ē���/�:��LRKD�DH�֖╾"��/�͹��3~hϴ,h���8o��-`�h�!�P��r�9	+:�	����-����{�����׳��6�����9��sZ$��n���K�ʱ|Rex:�X=VUK���Jƾ:K5�M�x��ڈ��u�5^b�x�;-��u�Z�|X��8�&��{c�bN�A����M:v��O�׏�S����	�+��n��V�r�]B3��#S'X&5��K��F����5D���㈛����,�b���La�i3
N��U#>�����7��7i��Т��k��3V-�Ndؼ��Qnس/}��r3���XG�ڊ��Dv����L�s]ج"B�`#-?���A|C�Z��H	g��Dh�v��k���E�&����=SZD��^�?Ih?BTQ&MxB���Q���'�A�.Rʮ��?}k�ţY1H`���	�G��"������m�ӯ=��2Sog�Mze�	>Ɍ����c�.t���S�ìw�q�U$�{���o|
��=A��3�v��0�� ��ނY�c�������.�&6}VJ�+���'At�
�2d��}g �N@$�0m��~}B�c�WW�O��R2��>spm���W��5K�!Q�4{3?��t��o@Q�nc��Zh�5��u�<��o���F%��rw���L��$cYH"����J��g *]5��6��ұ&�y{Q�vi����sw�p��q��,=�s4�H�e|���-(?7H�F��u,ms��0������ȂeW�#ֳ�߳��j\���%�9��[g�Fؽ)=">��t��w����0�9���},0����B�3R�T�uߖE�#�hrsǑ�%��f>�Gww���5�p3ݴ����}Y�doI/�J%% W~�o��.8��.���ۜ��0��"ȩ���{]h;F��T�.q��b@Pt�V����:8��཈�t��dj�v�F�P�%_�ɋb�!C"FG��ꃐ�;��E0>�#�8��6x�*�/���M�3�J8/C�Qߋ�B�(#F���;�s�*�u�vV\��3�N���Q�v�f�zv��U���0$��rB@�k>����qH��4-**[����pcݍ�	&��۶��F��ݚ!��|*�"��ߗ:��p��ro��{)�,��Tz����o��J��z��Ox�;�}!6���pTE8�+�&ytN)A\V�J�I?�a 吾��$mRN0�H9�]���kkG2��8
��F��;�X>��Q�hDZ7p ��X4*Q��)�z���ց�7e��x����G�h�����Ci��WW�_�Ņ1��$�Tz���Q���M�i#z�$�B�r�ո���:��9qG�����.��m�N��һ#����ĝ�6E����I=�L�T*�vl���OD&٪�%���ĜS0�;y�W��K�1�
RJ$�;E�2S����N��6�"
� ��ܹR������W����0=ǽH��"���|���4߂�D�N�D���US�A�r+�����M�-<2�Jg��E�E���y�,tb%"�Yw�x �a�ڂ�ipze���(gg]A �d�
~��ϢR�.J���'�C��f��G�K[�Z0��Y���f��N`�oq�7����u��.��	S��խ����ּ�ﶈ�����Tӈ��?;Z�mo'�ss|�/4�5�2V?<���N�t	����2���BI{��D�Q�?��IM��֢���2���x��`�<���L��}K΅��sRP�dB��؀�&� ?ʗ���9D�L�W�ҙ��Fd�nRL~�����BXt)�b�îj�6ڞR� 
��e.0^��ӕ���f/��v��{3�����Y�SaR��DX"V11Z��G�o�n�!GaU4���!b�* "�-�.~��0IyP�k��^��0��>5+����/�ɲo�����I�3��8l}SP�����^$�Mɥ��Ҡ'G�:�1���ǁ��RY�u��PHcWJO!��S(S  x~=|�)��=Z�M�����M�偦�G� �Пð��츧>~
$��J\���F�u+Z������ [Z��a�?������������B�,jg���,�C�3)~�ހ�ʚ���u���0!pkg�`��zFQ�)p���x���F*-	W��@��� ��_Ҙ������e�1��2&�]D���]t�����e��z��3Y�H���ٛP,v�f-�$K��_����βI�U�Bu%hJDJ��s�eYZ@�����Y���4s��8i������}5�d�`&r���	�����!3>�<��ˇS������%���(6:��
��?g�g����y�x��T%X
��R�zgc�Lf6E����|�������I�T����K�S�g�]���)��Q Z�u�+���#5�xG@g�����	Ҧ����8�G�#�?����_�\j0�\=�Ñ��YPc���-�Y���DH_Q�y��*�Iw�>Ƌ�(����1�;�E{�܅�'u�7½���">����"�[�(��؄;ae;�eû �?���c}���#[���� O�s����ԕ�3�A<�[��/�;]зR�sf[�-L�X~��'~�&1M$�6tU�ۈ]��ܬ�I@OB�_�Nj�����\A8@U��#ww�J;�T~�
E�����at0AVsvf����Ǥ��i�G���>|	5��b6��B�����nܕs�و}��=����U-�VB�؃	C�������s�Y��.�]���d���z����C�+K���c�]k$��*E��,l�XO	u�M�v��Ӧ/�+�0�=�ժ�t���6}	ߎ�8�G�	��͡�� �)�V
`�Z�o��Ѻ�G(��:��M��r��"�C��X�@�\4��q�2 �k�'�l�h9�1'�D>*�xYr�|";"�[���V��9z����ϝЩ�{���H�ʅ�bWvM�A"�.xAR��ؤ*o����iS�p�U]X��=<�H#���� �T�cU}��nFn�u�AoU��@D�[^�nf�:h�YU�­�d�Q�o��M��X��\wZ�ǎhU�	(�����h����ey��1HwTy2�Fb.Y+#���F��X�s��Wc��Fl*X����Z?�X�n޿k��n��i�����
�A*����D� ����X��}10� -&5�%M+ԫ�C�ST1X����2��Hl�;:�L��V([�����p����kd��B�Ez�!Sq�F�N��:�-�P��`�b����DɘvR ��D\��)f��=S��� {+=sm�^L�f+�5ϴ'�����φ�Y�[�(D.�����0�k�qΑ��o~[ ��E�y�-���t4☢L�C[y�S��]s�߽�s�q1yA�lL>&��:�CB3�G�(�����e0A-���8��Z�~�����A7?>�5r�5����'t����<��Zl��1��ɥq�>�g�J1���/��<�C�z,����C]���;z�8ͩ�,���j�?Ɖ($3� 2@ hWݥz0��T2+��S�������r�vg��3&���F� �b�l�Y�m?��b��q���)�_Z2A�'�C=lĪ�d��j� �#�1�Mwv�ؽ��ݵ��
.&q���4@C�,�T^��@j��(e\b���va�TV���S�����\�jQ.��}��z��
^>,���7��q�Z��9�1zd�	�EN5^>3��d���\ι\�����oP�)��/ᒥx�&��7�|�<,��h���؂�N�������:�D`�K%mo۵���{���){�p���и��h�/&����R��$yD���{s�s>�Ox8є+.&��GqΆ+�Q"L���'��qώjfq(�~b)�Ɏ�ʼ_
>�L�Ѯ ��N]��{��-��e-�0��������RK��7��3���Z�iNTlQ:�U�S��-��z�5�]3��]ő}�#^�iI��c3a_���v��)��2�txP���τ7iB�i�L��bM^$�:�?l5�����\!"�h6Ⰷ����rb�A� V G�ay�;P��R&�������ї0o3�"5�1eg�54[�h��F\��۶�w n�A�
��!�H.!�l̃�K<���m��]�?�J�ҴW(�2�P�ޘ�sY��[8Хl��Y��vi�6$���[�l����9�CK�=E����ҝ�5wh����2ض����J��o�},(oYg�z����|�ew��P�x�Y9"�H�ɾ�ʫ,C(M؝$�6\����|��s��:.Mч�Iㆂ �T�4v\yS�����Pn���Ҽ�\��9<�:z�:�H]I��ح��jؗ���_�ӯ����&
��2$:�VJ�-r��ݡ��Ep��v���T_�#�>OU�5�����ow�^��|ω���k��>B�D�v/ CDv�Y ��D�~F��V��p���8]M�~������[kD4���BB��ꊞ̶?�c"���������tH,�N.^��M�; [?T�\�j0p��8�N?�C�,[�P_\��oR�$�36]��Di8A �@�d̬�9��t��,�����^���gkx�&8LE���&O�i�l8��T���5�H��k|��im�VC�*�gX+0y�q�.ɿ�A��o8;��ϨJV�xVi�f���jS�%���}q`�תJ0�P@sbL���+J���h��J8R�`�/���5Y�;��s+�q~���Y�u��ԯ���Ӕ<s� �O~f���<ENJ�{6s���9 ?�#�\
j�W��0<?% _��ּ�+�����nܞ��߇����z���x ���
2���g	��X��vK�jo�-�P�*��D>x~\D��Q��nS��&�ύZ���ќ��!lB7գ�2�jS4(��`"{��9;�'�}U�)�� ��ؼϻ��_�?��������6���O�i#\�b�P��q������Kf���Ҫ��ݡ�QK>��B�-��������P�'ǭ>S�������_VT%��}0�SfYx]�J���~K��"XU�1hy&����l���3/��H���מH�L��X2S��6�KS�g"�롌s�R,r�
��l4��g9r����0��Hb�ö4�D���1ҥ��Z�K-	bf�[&�U��7zItkf-��HH��4�XjX�K�n�#g-�c� ���46�	Dt�Kl�ځJ=ՠ8����!ug<sBf�?č���ʹ�2��hZ��!k�PDgQ1��VL�[&D����ΐ��(��b�5�����;'�	[�H����	���'fq����
�ꎌ*�z� /�6/���W`��-�|����{�S��5J҆�sڧ'uo���h�Gt��R�]B�V$D	����T�3��c���Ks�o�1����\J�HAHM���9��⛃���(�)�E>ê���>:Zg���6��*���yYSWM'���}�ӾD��3+d��΅�{ґA% �*�|^�KDW��N^Jk5M�8�?��q_|t�ơ*W�E��2t�2?[��Z'�ͳ�:�:��$F0t��7F՞���Z�z^�v�q��$�XT��iz�/�u� 6S��TM|,9(DƼ���yh�MR䱙����s���?�.uI�F�w�����E�%c~���;�pJj���S ���MG@`��cl��K��j�Rg��l{팀?��'�j�Iט�w��M,ʔ0���%���J��`�oK,��I��}�
�f E�Ǡ����?�]
G���M�b��b��l�2���N~(���g&6��q���_[ƶ~+��x >֔'6a�Vt+)%��N�����o��]���oR�lQb��ٗ/�C`՜�Tt_�"��AQ�%��J�w)�W��Ip�h���8�5}Q��� ��!����=���W�A�������L�(r�#����S�,�A ������M ���0� 2"�ɏ ]��~w�.�T�s�����q�f��}󖥚�����7��ԞЭǿڕR@�%�n�:�m� `Ů� %�D2^#S��|\3����3�4s\�v+�����\����]S�z���r7�I��N@�	�VL�	�Vjկ��[!�jZv\�b���Y���\��>�z���~�W(̍O[^�j(x��s��F����[��,�Uσȕ����7p�x�l�&|(�� l���TY��!�YO�}�P��0#�gG�6B�a�(ٹ�Ū��fm�F=�ˤ�23V����]��;p�ʹ&��Fw�͉0�C�,"��a|���1�+Hb��|��w�YQ�F�>��8�P���cYiN�͖�s�c����h��B�D�1�Jv>[ Qu�zuR��T����B����S��*��ֽ]��ҿ ~���(���:��	{���+�D&�44n����
��O_1��J��Rݿ}pUI�N|-+v)�\����ի�&ⱮT������J�遽�RK��Q�����D�Nzsɒf���-B�`q�����"��y'��n~u�6�vM�)��f��:Fvmr�ۥ�r�'��տ�Ή��8��s^ё�,��Ί�A֑v�� ���Kb��[-yt��?�����U��_�r/��RgP;�� e�o��P���rk�z��84:?sH��_H����/���u��ٷ��\�`˃� Lp�����֭ܰ�)]�v�����R����?�q	i<�W�F�TH٫�ı�|J�l� v��Tn��I%N�h�2J/��l%�:w���y:�qa�n� l/3�ץJ�v��G,�����Ȱ���G��v����No��xu~�@�3�.m���*VS��P`��A#[�cx{"�4�;R����Nq�����~��Ƹ�߶�%�1��zq9��m�U�^Э�i�8Ұ�}2�m�	�˧d�Ru���k������Eʭf�����8�e����؋�ˊ�)�O���֟<JtNȱ4⁰����p#�cŗd�}��2��GO�u����,ucD,sO��쏭[
7��oG�(����=j�6i�<S�Ḅ[��B��8�(�6R����Y�>Z��J&�����YR5�.���W�==]؀<����>��XU����N,��Ҍs�H�SX=H����U�.c�?�
�D��T�R���4t����,�v䢈�x��B߰��.;��M�F����ʓ�X�ќ:�(Q��U7�^?Y��t�`b�"�:Q-y�0�/!��7x-?obd.�d�r�	x���]U@v������a�5#y��R�Sm�E�w-�TG��˦�d���ƕ�a���~Ê�Ek)�텺���V�E�p�,C?B)D.~��d9�=�sR hϐ?��?n@�}��@��2�_YϺX��-�MPf��	�`͜���p%qd��'	�a$#NB�K���.郢��x�lڿ�/6\�NEw�T�'촖�]5l!v{���j�7$5�OA�+�>m��y.Xj[��o��.�N��h��c�g���d�ݏD=�%T�y:��QDyz�s�+�d��6�rE�<�A�Q�]�&��z�Ks�D��?��2��4�}�g�g����f����J��,��ӂl�����r��F������P?9fP8��9N��R\H�(��fš�)Rq+8���ʫI��+�l�ܛ�����5TT ��(�E��G��Y[���1F3MMJ�;w1DB��8�x���=���­��fW#Y�g�3��9@ow����.ۛ����"���?#�T�{"�F��s��rG�Wڦh�x�.�ח��
[��y� <y<pX2�ׯ���N޹cG`4w�M���3I�HEYE�f�"]����Lĸӱ0cNm��1y�]Q�2�@n4���Q�맧�L�-�u*�4��'��눉GJ�$�d���'c�d˯�����^�xg�+�Q���D�:��	g�<W&��U(�bT�_i[���QRk���m�0J#�E�Q8$���x�j<�]XT\���6�܂�����uu��r��m�B�����ք��1
�ӕͶCÒ�Jo!� ��Ĝ0f8h��`�|�kx�,���P���#s�~`/\��b��yy���`^��8�5�4NzL�o��,�=o�N@O�`Τ��^e*����ը��l�u*ב�P�^�)Ѷ�sNt���X&�Q�]�<\T,�HR���ܳ���
�Z��1�v����Pؘ��3K�7��,>6
>��j�p��w��,���V�<U�3���+�](�!�����\�+��4�J?�"�v+q�NR�ml=M�0f����u��[���j��K$�[U�i|<��c��d�u`z|0����;gB`��s�~fQ�O8�[�<\T9�7Æ��_+���G@a)�kG~3H��}���& ���gLF5c\V��dmĈ
s�����|�N��5��͖V����߻�P��Q�&be��YZl�Q��Ƹ���s
E�*+y=�� �(�.$�N���u�hٛ�5�{�ʎ�2<��H�g��f}�ހ��8���Sao�=�!���Y!Q��M��Q@�6;9��Xy(��\~RƊ��l��� �z���y(۵:��ae��J2^'>c���
��oJ�b�6ìz6O�FbVC�tr��2�o�ժ�X���*}&]��V�\�}���� /����<��lק�t�vv�+RH	�z�8i���a�!qhxw��N���R����R6@�@B��<ZI4#��#�Yx*�?ַ�?�Һ#�����$&�4�F�%	$m"� ��{�x!���7�,�(kC	>�oX�N0=F���a�T�/��4U�H�rWֵ��>�"E�t�����F9�Q�z�6�\xRN���x>�]�9I��Y���(�Cw�r��+ܴBY9`�!�]�{ao��\$!����⡱;(:�OJ�3����%Ձ�2��RېxS<սw��)�݇X���G�_E���ɡq)���4F�dJ-5ݰ/-%\٫�q��znY��!��S
.����a��l~�;7xM����y]:x�C���o�z}~_�P|U�j��!�%��+r��>[��%'�L�u��S�� ��9EZ3�(s�R�O]�M��R/�����dp�A���
�	O�:*+�V_���&Y���ԁq�N��o3���I�{X��.v�&�8�<��d���j�%��̗�te�y�{��ި�.��tI�����ˣPL<�s-ŷ�Z�Q��!w3�䥥k|R��K���K�4���7��@)��ʮ�nUw�E��Kǖ�������$���q�Y�y���ͼ�#ǙK��� i"��pHݰ�c�R�Ԣ���'S�.a�iV���ϫ�[�/$�x1yi����
��3�N���P�〚�`���#Q��kv<X*Z��O�w�8��[�z M�^<Ovi�5t�8�8�ݲ��m���.C/�@�eVM�4Zӽ�ϡ��SFH�Ee��^��gg���d�x���DN))}�:��P��W�f���/���H�2@1�|�	΅(����A\��*�:׮QL#�k8�	;^n3�w# �߱�t�#Sh~G�#�,��#X��A7|��.�~�dbj2�(�-�����1�WGz}DnA��Kd0<'E�7��0�r9�Ҟ!a��-ξ>1���"�o�����ڹ$��N�����Zڸ��*��#Z~���=����v)�]H�	�'��fʲ\ꜼR����-B��홪e-*�ݥF��	x��J_���j]Q��JU��>5<f�K����]��m��g��	�
,��u+q;˺(����lGDK�Q�5�hn���Y�`�cOf�Ȃ�+�z@�(�#�nSt���|"`��`*@�|��.����[���R�/�)z	s�M��� ;R�u�z�f�������Me�i�G+���������?�M��#r��`c3�[��5{I�C��$7_�5Q��������G����)��1u���[��>j�@۝��ֳ��q����{�2�\�Hx�[|��0��E��e�����5���s�B){OlR�����Ţ</7�>/��4�m��e����|{�"+&]a���M����,\���I�mFc��d�g<Kf���>>o��#�Jڻő�o)��e}�8�V������U�H�OG���h��,�+��+к�,ǃ��w�۪%�^�Nօ:�߭k��mQ��8-J�vj/�h��(��n޿��z;9��IY@}�%�JB�>|�V�%"�6�;x���!���]t��}mp�i>%H��� �ϭ��ŧ���L���6�� ���[� u�Ax��'1s��IT'5Ǆ[�3�_أ��Cn�+��i��Ne��F�`KC��P�*�?�Y��W�d}{��Ư|/�zX�ʔ͟\������C�a�̳��B��u���dUZ��ްH�T���>�`
uk�7��{���1LAF�^��j�,1��E�{�n����V1�z��+4�d^?12��aU|�Hm�&���fk��Yr�,=�zP�Z���Q8��A����3�<r��u�p�S��)1�wm��Zy�k�)�yH�i"�HN����/B�ft�����35�I	��2~_���3� (�o5�,�~y `�|����`���VX�)�-�Ab�����F3���ቒu���kW�eD��G�F�B�<�w8O�����.˛����*�,�L�]6h�E��r�l�UJ�������%F�tW�L��ǔG��'rn���}��������
}��,���Q��Ֆ��e��I9C�4�	�L����$_�d_� ��^+^�,���raoY�? Њ��7�@��~e�����]�Rw��2w'Q)�]h�/���5�U��CUA��!d��_��Ʌq,Y��~�V �%
�E��r;����Q'�{j���l��;x��{i���q"5�l�[�N 4���K�r"3j��Ђ��Q�izz�x,��ƒ��K�����8"��j�U���&�F�C]���;U��(+E���y�B1æ�������S����B��h?ƥ�i��t<��j��u�g���;�| �vF��tPt��⎏ �6��O��ǽ�_].9�����7L )�,��g�@��oP� �*_!���-㙒JH����RD�"|
�GiM�!F��QdX:�O�\�lK����G"#`(��0|��P��E_����b��]�}�\1�B�=�?R�{����[�X�:oud�I�
7����ܼʊi�>��c޿"��}[���臃v"��$jR=�|!���E$)g]�o��-�埾<!v���?�����cWXD���[q'ԭM�m���YPs��P��ĉ,?{���Y!��k�ǭd	������AO��0q	�Ak�Q4��a���|��وiO|�j����qb�B��T�1��ע�)�dɥ�4o���"�i1��l�G��#��B��I<2Iq�b���l ��Y<�-�u$������yYG��̸c���YG ��u�%��;�i'����Έ��\�]�P�VU}�S&a����+�o- �~���%
��0�c�{O�'�W�pbx��ʹ&
���V��K~��uL�k����]%m�/��'Á��o̝�jY�D�����ٍ�EHO�j�[ ���	��x�g �$���|Hc�q3kN,@d,�S�H��u�\��ib�o�n�1�9���D)�����!�(\��&�^�]����$�9:~�tz/�,��'G`q� �4�
��̷
�">�1&� �"Y&i�=ci2Gn�R\��@`l���>�'<,�e3��n1����y���mnj��>�בK�;
',�<�ѡC���.�F��Z��j*��s�N�Yl�/^���[�_+

�D?����tݜ���[ְ�1?qYjB����R�j�կ�*6�"���w�}h��/�"��<�io�Q���;�jK�}���f��VIx~NW�,
Óי(��Yh��X`<p� )bb�;�+iU��>�+E�؅��9�U�Xna�T)̰V��9S�K?�spl����H�؊��/���$|
l�!B����q��Q]�#�+R��K�|���iWb���\%�4���N#x�C��3p�b�*���~���Zn��>p��p�m���^��(�~b�}G��U4Lxt$���FP�g��b�^""�c�)��
.]g�8t����A߻�%����n)�ݳ{IYܷ�Z��P���93�3I�u�a������fQj/���	^������v�v31s[����K��sU
�u>݄��/7��fa��m�za���Ь-�A;h@�8�5���40Ң���ŕӌ�H<`�4V�Z�^��%e�H)gM�[N�6f&���	���Q�&GM�1S��R�*����l\��hfmE�J�I��4򭰺%q�B0��a�<Nn�=��<nd�OOD7�]y,�h|�۾�N4�xPF�tU�z�-���!�Tk�2M'�@w#�p�:��
7����=�
��sk]\�O~�>��QtjS1}�&'W�V�er�H�Ie�"��w���Ct�`��w���n�.�Y�XUb��5b��=��ggi%i��d��_�����B�/fIE�����j�����]EЊ�9�Fi������%�$����!x�vrx��Sd�e���$��	�0GQ�@\Y�]f�hK��do)� ��~��>����eX�,A���(�I�m����'�{��N���1h���ͳfg���ٴѤ�w��%�~0@�u�m���++�B��!ڜ{v�O3y<���T�W���e5=Ó����d'�p�G�m=dU���a���!�*bL�\`�^`��K�d^ cB�[W[�������K�)+�f[^iۂ�
��t��0,�o(��^�o�
C�`L�o��7�ʏ�Ԇ��*��D�)N�Y�C�|x���^%�8��*~��(��59�|�l/,��y�ۦ�߇E��pZZp���Uɟ%V|���!�¢���w�eJ�^0(>l�y<�4��Ȍ1�_��ѻ*$4�=�Je#)p���%.W5���Y�摡KA3�H���D�ͥ$�~�� txQIr��Ktƍ��㹵:d�C�V�&�mn�dH��c̳ R�{Q��+����j��^#!�la��0�dͰP��_&�‾Ek����o�wP����7�ʁs���]�˿9L
�"�o������ƻp�a&��1����!�pp���	aw4�0f��EG=ih�F!��q G���l��0'�>�(#��ҙ{;��Q^i̜~���7���\i��h��F	>�W��b���<:8��+�w^��+`��y6nn:U�꒥���-Rۀlڤ ��7d#�dEd�����7�iX���;�7���כ��Ǫ�OJ��#��a����$ *��~��pCۡ5���>�R�E�^,H�S&����>F/�7J��&��=�:�|��>9O���q��ƻ�ͶTI�o����1����i��Mh���5[�ꊫ�Vu��|z��ń�pU�{�k��R͏1�&���̟�	 ������w+O>C-�FJ0ꓹ�h
��}S��r���!���Y�`�NH���΅���`�_�Ţ�	�5��2��FMN �VV��	��L�.L� yУ�TK/�"'��L
P�+-��=U ��=p����u�7ˇ�|������n:=�b���뮖s���o��{vJ��k��>�.�|�W�0BnU�o99J���z(��w%���P�}U�C�������_K�|`��w�R��oX���dϦHDO�����(N.4��b"<wf:�*h����l�0�?��%<�����P��ol�����g�ZO�C%��@K�����N�`^����xL�V���A�3��Ğ�Z�i,*�-��l0mߌ�9Ӕ�܄}nQ\w+ޙѪY~���֣�P'P�.��0�Z�ﱫ~m�Gjl�[o��7�_��N+��K��?����X��j��ˁۤj����_'���ָPx!�z)K>9�N� U��H�؎�%��g��w	�AEѡ#�n*�Y^�$��m0��ې#N1�L����U��v0��,^��`;YI�u�؄<YWD�U��q�� 9PۣJ�����|.ݴX[��g�ӌs���۝��� ���6ԭ�҃��.I�Aխ4Q�7�~o��#�7��h�Ja��¬�M,�j�Tg��!'�Ob�/vڱ�Y���U�ة:W�����Q��Gr�x�Va�$��}�����ֈ�E ��Z������)p�Rb��2A�Md��U=A��M�c��W���}=�M
�~ɔ�R�K�bC#�^�,���<ª/5u����ף��@'�@��ձ�.�Z�%vז����Ȩ��>��WK7f���"̈�c'�.��G�Lr;8
ϳ>��(��x�߿=�o
�Lcg�x/�Q�WOj���ř�O� �,4�~%v{��8�]Z�y�?e��W���.<XͰ�)�#3B��x�Q
V2ƩS� @>�\����B�hS���]�I��I	3��P&��+�L@�F۫k����(�:�d����3荦��.t.�ޒ/�No�~�訜S����7s1��8\ƤԶ�V���DK�h�xG�׸a�H�b��g�s;�sf�����o�%-�d��F��?�x4�t�C�C��m�|�˺��?^�kkщh�<�h?
�[�Y�搃<rN��X�<�U,y�:����rt��5v��2�=��]KNY� s[Ŏ���ڏ�{t,��`|?G���_a�+3�F�8/<�9�Ǟ3u4�Ͼ~�|��"~��}	P���	�s����x���tE���$�T��:2&����C���=R��d�DTf��]�]�Rٞ��q��.v�BL��W��aL���
8m��w^NL�xW��7��������\S�%u�?kI>}��t��vo ��{��®�c����*��N7��4�\k�G��Wect��K�G�/�0�B�_��lȠV~O�
�zy���3�b��#��do�B��`�@� j�J+�ؽ���������	�I�GwH�;鹉�̺/$E�f"lV2}F�ѐ&�g��) )��n��EO)E��Bc��6�Mm�;�1 �1��(�%��O����m����̙�%"o�{���O;�����#^?�^Ζc:��(���i(.�㎑��Z~(ێ���i��[�Ya�!vT������:
�]4��ꭁ�9h�d}��/��$">B��].-��Yi�roõj);�<��i�	�Jce���:���(�����40�#U�M��C�"����5c�@����P3��-.�_ >�}m�����G��tb�����,XSR9���%2_S(A��ڴ/V���.3�n2�6R[�	)�^��@T�j���#�(�g��:�bQ�;v0����o�ı�$���� �	��j�u���-k���;>P}�=�����%�+�P���V�z�Z;��x�%�Oҙ�#if+�B:��Vvp��>ӓU	�S�tC0��~>	��U�ۣ$In��z�yPI/�θ^�P�|��$˽��jJ�ΡP1l�{��`�3��g�
(��sǖj�J���CB�F���{�Mtӟsq4 ٓ�y����:�C	����:���1����h҂�Cau���O�x�g,���|�"�nv6$F�f*�Gw�I��Eo���&������o��)s� �`�<*h���{y=���J��z���"U R��Mw^q��;�?f\T�.�`"���YvnzgRx�o�?��5Lf�r�w�	�w�j��w���<	q�C���:z�־Ǳ{��W��N�H�hm��������w��h�9R�^T�y���˘[DI?r,�N'�nc΄��&�j��VY���[��r�M�w3���l�~�(�ɢ�)��Y�d@s�Mx����e�W�υ�fY��4�����%�l�^���T��=��`3z��4��&�-�u�2b��"&���o�W�HAB�����9�bظJx>tsNs��7Н��c����^��n��`����&�Z�[J�OG)�}�*�ک�u��PP6	E5����	�#���g�J���&T����]�������m[�Q��g��1�������\?��y+�(��7kp7U?����3c��Gu��T��-d��"�6�ӄ�p5K���g�T�oG���8H�V=>�㱲/��'�;�W����Z�m���.���\�H�F�*�jqa�3�>�9Z����	ܗ�t?1~����;1;��wٙ4�o�V쵱����=�]}�y�b.���. r~�b�WiZHġ�݉U�h�ZQ�/���j��X_Ɓ��;w4���'O=W��Ք������*�%_{3�d>��|Њ�o$�1�Z��M�G/��L�e(����H'e��Յ�� ��K7w��Wʋ���`D7O�#&�8x�]�v$֗�Q5=�2��.�58�V���
Ģ��b��N|�����*!@!�ud]3��G���ḟ�V���� E�d�V��#|�֜�:/5����@=��\T?���:�p�!��:R��ԑ_�}�P1��5P�z�B~�z%,���'~�2�$����
��i&'1�w��{������Oll+�#���|!���f�O���d��
����Я�&	K�i���X�n���x�l��m�T�\�o���ьk����n4w,�����#6�w�~ʭ��UN�8�=lӆ��t��ڏ8���'u�>�B��-�o�vΔ]�ĥ��<�EĽ����I�,��2t��x���+�.�1W��R38��(�|���6���/��bW��1^߈7u�[�%3N�T�!H$S�3Ke��j���V�.T��R��(��ѿ������A�`L9�+>m ��oiQ�f\�`��؟�4N_���'y�lA"���2�$�ߩѽt�jѢ���V�X8�n��j�a�t����Iy�
/��W�+�`Λ�X*�|ObJ+��u��U�EjkIT+w���֟���G��*�����p����tW�t��Xq$�`b�R�'E*|�,��*2T���A�_���1_�6���H�e�WM![�l.d��mr��Td|�ď�Y���YiL���]����dU��J�/D��x���'=��
��Ԅ}a���� Yg茔���T,}M �h�`�Oa����7Y(U��6�h���Ra7���Ϛ�����L�e��_;M^��L-A!����dHt���i����b���
�74�r����F��s����!��,�l�?_R�}��	d�q�K�b��qD�Ë�\�۠�ő�L���>g`?�gg2�Rƪ���[۵�'$��P燓n��پ��^�Po�RX���Ȥ��"�X�b��g�(�̎��gu�QDv����P���<�<�}t���<���MAb�iV�)ɓ@!�C�[RL�!�l.p?-К��; ���;r*�	�~�Ҿ��}K��i�K9�[�|6@��J������k�1�����VX�=t��M�D(����L/�*u�Pb��p�|��LYu$2�7��_��WN�W$�2/�m��j��2ف��|5��7�1���\U�ju-���O��uZn�7��]�zzɘlD�1�4�t/�.+�T�	,.���Y�3���.�F���Q�yF�Ĉj|�({�*���X�����do� ��[�Żք��XG�F���I����x\kz5S,�>�'pT��?�0�0(@=h�Ay��Ԝ�HY�f\��DGIr�KC�V}�$Y��xn{�H�p�	ׯ[�F��Oݘe˘$EG����pAl��wSY.�|}�x+����;#��.�(�7^��n��ZaѲ�����D����KaH���KT.:��0k-k`�l�NO��݈������� 0`I�G"1�F�˟#�ROv*��Ce	���)[�p.��$xH��Z�> A^a�|v���Mr��S$�_m�Qy�$��e�^�i�v�4Xw��v�������.��YL�YX�Y�ب�vNJ��NQFH�ˈ'�		��l��J����~���
�s��O��׫oo�{�����(d��2��C��M�}ɡ��1��6y���.�rv�BDj�8D� Qx%O���ְ'���fA����4��!UD��?K7��
��ܛ#�r�;�bf�R��Hr���JAڏ_�`0R�1 �B{`�km�n�-��wcⅽ��>����/η�p�V9�䭇��!���+|��#���M�f{���'�4�Q�wZ"�lѵ�u�p��N22�	@�c�� �����q�!(dS������i=f��
�� N�>|C�$meh�Xq(S�C_"���X�Xv	 ����ǭ�v�ǌ"|���O�V�O��vۑ�#`a����p.��/��$VyU ���2�0�{/�Yg�qaSx���~���!�>�~�z��EȀ��(�[o���<����q���g�ܢR�`ޑA'4��?=����`'�[��k��\����� z-d�Q�_�"Lna������9g�oằG�ܖ����J����pch��[���Oh�IV��rcE���0��Pc���C:�'T���_�X&v������T�x킟�{Y�;����ސ��z1�>����.�.������3��>{;����6�1�k���|���
��"Ö�Q`�NuM��s
�XP� ]����&���#C�ǚ��i`|oI�f�I���ev�q��^E�H�" #�&B�C�;z3-K�Mz�P���d͈&��/�e�׺�>ړ-�ʉ�6�o���M²T�'�5ұ��U���nfUfؚ������ўY#�����Xb�#���r�@���z7�JB��u?+Yi	����,1IǗ�5�/��m�/ ���s��x��B�4;��\>T��p��׶ƠD��*�8^bkD���$o]�\�+�jNr-��o�лݚG�a>ب���[�"�%��)Zf���?u���[�0-�T��@@��(��`KL�V��_MIg54]�l�g���@�K�B��4C�E���+�9�ʰ�~,<bf$!�.yv;��:ŀ��w�c�#�V�(�u�N�h��;t\\�GJo�1�<-c�ü?�^��;K�O(��s��8Tv �*�(-6	��v��eʸ\0Z_��4�	�,�b��D���&.ib���fQc�r��MC ��w�X�	Ɣ&��������3�i-��I��'�_�+;���S|K�f�|�g+�}��C��S]�w38棇��Ƴ�-�F�c�=G����`�}��&�!f�S¥-N����5�ۯ���T6S�M#D��PSΫ�1�,8��&=������CE����+9���5M���D��-�����*XꞙT��V關1FH0l�""��Ғ]�oŶ����ul�o$����g4e0`}�Q'jA�I�Һ��\�+dC�<ʟ1>��R�ж*J�D?k����R�Iz�CֽҸ��������A������:�U�!����R.�֘*Cu���<���E���p�MQ�m��\�P ���
"#���#.���'!j1�3�9ϯ��(~ͲAВ��� ����]�3s��ŀ�JC���~\%3�Z�}�Z��������"zΉ�ؐ�# &�uD���R;����U��eր�J�����V���X���%�f�xx�:�#6h!�W�6����Ӏ�{0?�6��ci�\�����>3�4q�$]�"$�7}�䕀B�vv�P����jM�XH����=�tp�h{�V��,���ñh�Y�Xښ3�r�#mް����zHވhB`�*\�O��$�w�	ʾ����ܷ�d�fR��R��FL��ކ--�84�r[4�2���%$���A��
J{m�Έ�D�(cJiEtё/�i��"ȧ)n(� ]��R��B�<DK�* ���]����Zm�/����0�Z���yE����a��I(+�G�<�V� o��1�y&sA� �lχ�K+4�_%}�|ӡ�MFv9'���`��Ɇk���-$WnI.t��4Z`��_�D����Q!�@0l����}�~�ct����V���?�Zu^:+A [iNv"�éL�O�ꁣ�:�xB�p^*׾��_��G>� �O@}�J-לd����Ey��l���ᳵ��u�D�>e	�{�:���B����tY��d��uɹ���{C�t�&M7���}WC{�5���X���
���-�5��=���)��X�N���d��)f		ѰVNir(^E<O����v�*<�`�e��IR*�Ȃm�Bq��$���Ɛ��eȪ�>�#L�(!��*0��9�t/�.��ym#<;�"��lT����R�2����7wf*n���@ �$)�)��2��ؽ�P-t�zk���\�,p	��t^��Y6]2���{��%r�3!&��bX���l��]�6�`5��I>��ʯ?�&ɥ��$��V[]s5sFV��'��ʪ���{<8�=�/|�M\�
(��@b��`����?�b�B:={�b_A��(�$�I3㔴a҆�{J��T��I\�C{2j����*߁m�KZ�OkaoO��/(�,���M_�X�L?���7>e�iUb�(2��r.c�8չ�*j�))ٲ�|7��9}f���-�=�~�b|��3�˔a����ˉ�R���]�&�{����X��i�笗v�������_ �J�/d��}�Wv�E)>b2ڐ�Z.S��o@%��q�ݕ����sQ�eɹ���:p�s����5s�1���"��D��Fjh��^�����o]��ä�E*p��~�w��\��ۭ./%R݌Q#W�'8X�n��䖺�~8ݩ�W�խגDo�*��uJ�d�xi�T��B'�D���?^�#3��S��
)�e�4��r�į(��DJ����$K��kRǗKg��V}��FK���ǣ�(��Y ����Fy�>m�n���4�s�Z���Ƚ�	��ZoG�5�6��9.��d�.}�U��ͬ��?�=�T�C-��u�m��I�+'4��n؉��c��e���E:ZZt^���.��z�Ի6ԡ=�����4jU"����,n*$�h���;H�Hd�Ѝ�3*���� ���	T@AĜ�������;�A���֍3�0��uF�O����mٱ{�(���-�Z��_��~9F�d�df����J��M���鋶��mT�H?� ���������SvE�� ��j̮P\n��U=}�hL��<�9���,��#�ǆa�5y��3��M�S�����E�7�c/�>A�7��H���jl+���7!@Fn�܌#��;��Tg�{Q��&YI��Y?ZO�W+�َ�f��wL����u�$�O�P�	�6��ɳ������_�o�������~��82<L������ɌTu��>|KK��K���!��Һ�e^�c��0��(���U.\A�6ꝧ��O���� ����<kƍ��*�jl��B+)OO)�&9�:$�!�~�qw1fyi���)�,D���������m~���?%�-��;m׋�k��>�xInMt%�ǍrS��D������Y`���CF�\ ���t��2Q!ȝ�k<�IOe#�}��R�2�!$���zB,�A���㰓뺲~4����1�zH���C8j� P�P�Y:f��P�Z}�;�#�)O��<._w5J�q��Lg�rJߏ�Jw�c����"�y#`����ih���}{`����m�@�)�	)䊇N���?uI5�g�'�䁺����kך����+%2�A᧷���/�q%k\��fbdY�P^�T���������
�J���/JO���W��c2�j��4ij��̈́�����(h{��z'����lRs�}Qh�97a��nl�b�~j�����b�n�?] ��e[v�K����k=+B8E���b��E��%�G�~1��kW�]y]����(a��O	�{?�y����W7�Yfͨ8c�A�����e����tȍu`s��| 茬sg����Z{pH}3���*,��BY�1�V�{��S<pǧ�~���cKZ�Q�f2U	Bwg0&(��eL%�Y�	}�����x�y��A�$����h�O����4�DT�/����Դ ����u�����h��P ���yz�==��O&N�P(�;$�g_�&��;G��j$�S.c*��ъ�7�p�O�,�12���ԑ���PI�K%��[��,�-�oOa4�1�6�Ay����x��`m��v-0�0zȮ�Kv�̚*�V*�wa�YUM��oo�_4MQQ��Y�rGnT�po�`��%�f�)�@� ����W��S���SA,*�v��ڈ�|z�nU����#^�Η���P7pMt���)QQ'���#�˔�̔-�{��&�_�KDp�sY�dB�B?,��%�j9q��1g�M�O��@P��b��i��T�Ҽ'3��Ѹaj$�ig��ؤ��nK��z	
6��"���͑�D���:�*�Q�� �a�h��ז;�&�:�+N�3Ɣ��P�@kl�R���I�8����U:]�$�a�m7�T��w�a��ɽV��]��|t��9Ϊ���~/�3<Ƕ?�,��a%'�7I��|�%B����q�<7������@9&���Vqr��w�6�F_���_Z~Ղ��;F�KM�h*8��p�s !��{	m�&�y�/�A�gn��;���V��"�*�3�����3˽�������9��J�3�;��Dj>W���<}�SY��1ۍr2��j�|4��n8��>N؍�ԧr�7�ed+���;[B�SAn&+{��*���{�l���9O�N�������K$�+�W�׻k���jGr�k;�S�[m�KHa����ו;V�&��@�/F�/U'0�.�g^���V���hm�`)7�<vp�I�#�S��U�҉���3��Z��F��I�=0�zLS�?ͭ�q��F�4�I�Q��ab(�e�~J]�}F�t��0�O�U[њ��,u���Q���0T���D�f�S�n��k�^����<��6�({b��bI
��@[٣" ��0��xh4�ʸԏ_G�I����>g[(G��2'zPqA^E�OO�g�4a�Zg�s<s������_��F�Oa�o*�{
�p��J2꭫�t��i�%<�����Gs52�}�h�B$�׬�&��*?�
�p�l�]�S:6!�H��P������fP�&�_�ۈ,.To�ֵ!���a�o3�B�Z+UgڵW~��jU.�P�e:��!B���"��R����V�c1Lۏ�o�,�{���%ic�tw�	G�c�$#E���7�$���t�au;��Dl9��˅a%E����^�*�B��@��oO�3+|\�n8%��0�J]�3_���9�j(�;��b�Җ��p��Pm��!I�2mM�6��[y�e��N9ٜ����,�ஞ4;��˽�Bޜ�)�"]��S$��큾�u�����c9�hVGX�Ɠ�[��|�]*�O�@�E��zèC�{�S#cd��CI��[��	�R��&���FwŴ����[S{F�c��S�{�4��8Rرy����|�,�қL�a7��g�6íJ~�	p�6�(-�sBߞ�Y�!�~"�<?:L�Bs�;jW،(�X��t�eKLO�c�8ig��j�  ��l�H]�NF�h��@ e^C�$49����3u	ן}]��R�=�����}��D��V2��ǌ�O�킭�B�7ܠM���pp�Ǹnde�7/�U�C����:0��S�p$�Q M��4��{LU��Y�w�ż:b���V��iۊHb��Җ�0R�ۦ�%R�L�F�*[��qC.�+��Gq=�|~_]�x���w�xa�6�^WOH�9y�t� �@pw���M�
5)�Z��&U ]�Z��=G8Եh��<Z���\q�����9~�hm���B��_����J	��Srje�?ָ�S�ܨ#�?�OOd�_8?ʮ2ֱ�x��q�O%`��.eq���%��F���9E�<6�4�,�ۃڤ8�7��&EBv5<��u���8CZ?�.V��8)׾z7)x�U?�=+�ڟ�لr��V��Rf�,4���d� .��RQ5�\��������m&�gL5`��i�"�m��lؔGQ��������N�+K\{i'KhWf�Q[���G�B�1)��ӗ��|*�CF�y���rY}ₛc?TM��g�2���Ф�M��:79�l߇���7����H(�l��'U[G�[(����� ��z�si-f�+��R�5��Z�A�2eS�`����ވ;�	wNf"�R��m�g�V�<��3}�lL.9��ڎ�O���DG�Nk{�0fru�&�A�6��sM%�g�a��:����''���p+%R�lk�&%T[��c����Њ�\�P����ޟf8|{]��}��ӣлS�����‧�o��a��@�}�i!�!i+��H.7>��k;j�"��R�f��t L�p�B���S�ז��N�!T����'\x�J��r�,r�࣋�*�~N�����.�7�!d��XunVx��;�	�R[rs��j������2#=����\��"�d���sT��ְ��P��
n|d�^��I��Bےm�w�
|ǿ�:%E6�9�������� `���w������ؾ�L@��ڠ\�c;i�Q>�S�x�9,V�y�H�nN |M{��^a�RX���j��x���&����}nq�>҅�������BިV�\�tT�v;3����L�ƨY��t㇊��|s��ޒ5�����5��������;d.@�/��"r�p�Y���݁���D���s5��2$��Y��Z�3ε>jX'
=�	�N甩^O���ޏ�bl���1
�:N}�0I�W<�Ga�"�?!�6O�%k�xww[$�P!2���DFFg��j�_��d4���%�S�(��k-�w/��Μ۾�v&-/������2N��f1X��=�\&[pF��Eg�K�˜�Eד�^S�%,����M���T�&�d�;%�d�(���}�X�o}v�6����nfS3pH��@�ENĭW6u���|�����[���㍍�(b.�[q"L�Y��*�~گq�^t�Z/�z��@|�ދ��JÅ��Lg�#�I��-����f+�i�я�(���;��^�e���ˣa���dxM5޾L��m���[�1����*DL�w�[
���J�TB�Bi�~�?_������i���\ަ�έ+D���>���ط|a�D�wI΀��F�K�t�����p�}�fc�xMQk�ߊlT2�-I_�zW��"h�d����z�����J�$�l�NP����D�S��[��DK�1M��f0��<� �B l�k}"f5�6���ZvP~�����_��R0D#�#u���651�enzA��c/��F^zDI�Z�!hr�\W2C�i�L�(�CJܪ]�p����H�f��:�[Р?�d���]P�bA2�_�+}X�^k�.-ՆZ�Gh�^�{�e�� ۼ�(�(ܣ�nty��F?�ݵ���Jk�gv�U9�nO���>q�G�{��{����d"���]S�Ͷ��g�`yȳ^WM:y�(�C����c��� ���%�'d�����[*P�>߈^C�g�o���Xu�������]��ٺ� ����=١�o5���/�`��>���Ƈ���o�f�@1O~��W�P �"�OZ_��OKa�����_�`��D�hA9{e�M�	���|Ӝk@p�>��h��` ��=t������h�VX��g|1C�V� �ۀ.9(	���?�����_p)�y#A�~���%I�J���k?����A�>R��y�܊ca=H�䍉�P����7nn�{�*��
 ���ԤJ��3�m���b1��,�T5ʝ��A?H���������X-��B溂	b\��&ٝr�pP���o�u�,sbJ�z��jr3���I���ڪ7Ȩ��b�)�v��O�3Uń���;nO��\%�Zy�lƧ>M�]���=�Q7�A���G�cOd��#�ytR5�_�zȵ4�w|���j.Y�,�I���R����t�����!K-B��ω��O�˴ť�*����0	���53�Jެ֤CCF���ghz%��������������w̳��a*��a��
\c#5%��pT��X�o�<��ɋ��J���7��%�nP+!k���[:�9���i���1hf�if��Xn�a��A��%.���}`9�Mp�m ۾i,!̷��~�H� ,Ȥ�fpq��+��X��z�H��r���S��	$�@0�����(���M4Jk՗��V',K�$�Y�ԭ����4���N���>�Ǥ)e��{c�j�?��jdg����/�� ��"*�EmYC���m?7l��}����5{o>�[r�x/Y3f��9��w�I޺�1#6ʚw�t�.z�ey���ԥe|��ސn��@OHt%v8g&�a�dn������I/�(�iZ����YD�n �&r�/����#�\�QD�r|-��ZL:MR�\{2i04�*2��N�`Nw��W}��s^Ц�	-U�,�w�j�PJ�}�6�2QvV	*C���~�iRA\o�Rb�e��V|���o�~�b�g,��B���b�:,jf��΅0��hxV�(Ȓ�]�~n�&��Zb�f�GecxZ�,��X�M8v��N?��nEd�h]�z-+;=y�	"om8,[	Z,8�g�Ĺ����������q( pnh�^��7��.N��m�p���ƥ���E5�I��S.�KZ�vǠz�$����,���զ|呥��)��0�Y���=��&���ņǑ�0���x�~�R�C�)����?�\j���x;r'͜��D���:B`v��*8"�g�	�����#-��r��2�%p�H<6C[�ߟ�[YtW���.I��IH�'L	����ѢY%�otvs�����C|l��MEᩀM�44|߿�R�l�+Ͼ�'��h;B��A��Me�`�su5!�'nc�J�v��\�C��ZP���x*�y�wS!J]?��L��O�-�Ff,c��V=�{H��R��_M~`���)^��>���j�Y�I�y�����Mg�<K"V߁#X/����i���`]mъN��b
m����$����Y����g�I����YH}#J�3ع��Nܣ�*w�t�8�y �d1�ٌ hio����f���׽��I���J<�����l;P���y ���N���t��[<��ȐĽmm!JǺ]o�$0D	��L��n����[˦��1r��c�B���.>b%�آ[��SLX�.E�[F�w �1��x�p؅�C*�`4�G�`�s��5���D�8u�Dnt�� ���%J����'<�Q�:�� j�X�
@��Rr��&�#�x
!c85 �ij]�qx��T��X��y�O�sԡZ��yY���o>T�SZ������BOC����N�f�L��|���P���z\G�'��R��p1S����e�pЀ�,Q-X:�[�pA�O��3�o���:�A$��%yV�馫 E{�&g��c�Cp���x�ݧ2��S�z������m��$��CwV��YQ��P%7c���`��)̤\�$@���Op�K����L�m��_�|��6�I�)�$�|���<.�����wG���~!KH��D�~9o�c��-�o�ʊd�ǁH4y�����NЄ$��[����zh{u�I�L���-<��1q*���˽�~dTl�E�C��H�nX,(;n���=�3x�mxN�rL8�ӁɧO;W�#�B`S�u�ў�P��ڮ7��X�)�s"#Q�ĦT;b�߿/��0���..��~8)�]��WEZ�M���i_pc[(\+��ͫ�wt�������~���W
���ٛ��&��RAX�UD^/���nq�~�sy���Vt���k<@���i���;�͕��*�;<��?X�"�K���>��iц�opW"ɀ�v����&K�j�>͔��4�kB��k3p#7E�T b�EȽC�b2�R'����������?9J��J�趂���Ь.4�������6ba���Xa$�@�!	�M��`�f��c�om�\$��܆��(�;#���yQ	�pF�����0�X�vK�!,���k�W52�.�M�㭐���Ӆ?��Xu�Ǭ�Nj���x�ڏ�.ꢋk}�0`�MMrD蜭t"�d&V�Y�fS��7��%�щ�"��̴'���r~mř/����*#陊��\���Ȋwz�+���Z�f N�.5�]Mu��_���&��Y��O��~���v�,d6`���t����P������<sLQCt�dz!)[�O9qJW�P%�kdzp����c�n�6���2���^�>f��631-����f6��Չ_p�nD��ҡy5�'y�ʸ��ew���_r�h�K��M������������нu��m���SmS |��4���Ӝ�7��ۻ_^�'�]^شz�.	�<b��6�%N���<��Y�F��8���V�%�?���+58�(��iҖ_g��-W��`\D�*���	t���+�I�ߒ��M����S�ۚ�3p�4{MRo���M�}��#����@���Nޟ�,�"�=�&n�w����bزE��y������w�����۲��{���9����\�,,�pM�Հ��9n��w���������е��t��
J;��a��� v5b�V�꛸�>g3f�k�RM�8�`G�P��Q�-l�v]�%�*N�jbk�C*|�`���(���<�pl��4p��/�f��t��ݺϪMݿd��
�zF��3�0����D���]��#m��8�#���::�Y��,aV�R���K��7���oꧡZ ���˒Ӝ��V�;�Տ�ᎉ��& �ivh ��>i�{ۊ��ǔ���6��U�lQ5�QF��w���KZ,<=?���M��+R�A�����LB���u�⇤F���ڢ�=O�B��蹊^劖.o�]�����X�`��$\V�.�n^{��e�,��w��aP���J|���̇b[��!nu��i�6vP�<�t��E�(εg��� Bߤ�����8�I5�� [.����3ڧ�T�;�(DO'�z�Ë yt6s{Rs���~���
?�8�MK����������n������-Gg7g��l&#���X������A��� 0�:n/��94g�`�.ڌ��JXjg�;,0k��֊��v�fj ,bB�n܏J������-i�"�%����g��A@hd ����̎�+)o�f�N
;p%�O�Q����i�T@����%VY�:Y�Q��^F�H�B��0�*Q�:�G⁩��py`)B ʶgPW��	�yc�m���ӆ�K\�3�,m�
�p�ʤ�r�b��)�g��}��vN����E�D�Ň��ę^����m�ܥ1;��!�/����,�9�>�2����w�3�I,���]�?�l$�����2�{�oW´���C9h���*!46=-������9 ��� [X��8�3��5�i������>��H>��	��?tuE�D*�p_�ޓ�9%j9���.e+�o�"�g���<Q�p��;�a�b���9��5dd�?�O�,)�)*���M+5V�B(�5Z����ǻ���k�wq��,�Ui�>�9�9{�%/_Н�>1�X��$��V���8���]G�&W\�' kV���D^h5�3W2�� XK�2���.�b5{�4״\wK�z.�ui`[ԣ�.
��Y�P��ݦ��T�>�[��"_&�uR6�~�O��QDȈ����nJ�=m��ւ§��G*q�1#%Y]N�P)P9�Dӄ��b����S_�m_���԰(��qz�KD�Pf��2��,�j�G�S(��!����0�^�����OC���u�6��+��-�Bp7;�iNx�]�$Z�Z�D�� ����;"�y$�7`T����w}�k�m�0i��&����ek�w˩����&��C��?��*��k�˞T�w��Wwl��*)zĜ��q��9�s��b�0�֑ى�)��m�����A"�u���`ݼrt`z�@��~ͫ��gI؅=�֢�$����M%?�:�;�Pn�u��X� �wy�@u��]×Y5�I[�2ǆ2����(j���Qa.8iu�����sv%c9q��?�A��C^���$�������{t�����_����ÙA=5�-�#�6��;��]�VY�;R�֋�Tb��/��9�[���r��v��Y{T���(5�Tnl�*=��U������vC:��U�,&˅�|����e{-N&r�SXl9s>��]-4հϴ(��.���i�w��$g���'���$�O����O�3G�i�%��ڇ�p�dmN�2�]��)����yW��q���;�4۸�0�Y�)��i�ɍ=d[��fƞ.ܻ��Z��C�YR�^tL��L���N��s�vL���?4�^&͎T[t�d��<n�"Ru$���M_�_�c��yQAʹ�F�FnJ�IB]։r�:��
��,�u���4D�5�J��<,n~'��=�=�m�x��sF~����#��Ψ)��oe@�>͙ۛ�r*sF��d���	�:]C�B�� ��V@�ם�,�Y����J���������{�]��h.�Z�j5�D��'?*a ^-6$H@�A��:[�t��W���ĭƠ����%n	D�$^�+��n��H�o���︢�/Z��nd@�Q"螫�� �sw�SC�U7��)�C�]/�'���QY�[ �2�1��§^
�GX1=�z�7�c������>5ʀ�-`�� �I�3�2�t�J������.y�L���7,V޽t��J��QV�R{q�
p���R+
�2ǹB���p"M��.�-%C6fi�*��K��9߽�=5���4�=&�"�qc,$͎��R('�<Ķ(m@q����+�0^�`R�Ms����
�ۄ��%���:~W�@ݩ'K,)�y�q\yՁK�O�r�yiVu�?ۉS���_o�l�z�M@�/�:�� �q�g������� ޳usЦv�ލM�H�g��P��++�Ѡ�|��v��5�(�-9�Q�ρ``�,$��<&
z~�%��lmlfٰڙ}��g��b{�#{F���3�Ύ0/k�#ZW�����r/�S`y�F f�*�Uy�qV��7O��qh̹\�%� ���z�8ݍ-��i O���O<�F3�ƨ�P��ʊ �&+]�v4wjYO	E�����D��nj�F*kW�b�i�<�o���֩@1���0t���N�~1<$�h$���ơv'�F��5�[r^&@�{@�,!=�5�F+r�t�1L�ԋ(�|)���G�G��	ء�x�8{�(�[DN�7����)�v��,`�F���_R�k�,�S� W�0��-VT��אe����iH3��fq\�%PtZ�B�-��VΉ��8@�#�x�፨�������y��(_N�� ����6��T��)Ϫ���f���5�����[cЧ�� ��X���$]0��P�oO�y�QB���6�"�P�'�C�ψ1^Ibfټz7 !J\2���+��D,�K;%���=��8��p]���0N��ӲM���%�KBbM?�����m=C��@)A����^gt{Ne���c��>�?��$7k|�����}5C��I�`�p�[���"�A�V� �@���w��<���3Cx:����������B*���,|}�i��������
.��p��k� �0��?��������Vc0�|A���#���u�o`x �b���4oDԑ6��V@��Ϩz���~�ْN��Cj#1G҈^�n���=B!'jB Jc��M���	��	��1N�k>�o�_i�z����\�*�$̦��h��3d='~�1T�M�(��ƨ�]��ܮ<*��۱Q.}o�B�1�u5�sM�0�̬�*g��b����N�+;M���Z��1wN�^�$Z8È
R�V��h��Vk�X�Y���~�z���x�'r���آ?�fj�4��6�"� ���-��ڭڬ)SU�p�C����>�&=�D�6ص��M:�U�@^T��]�C�ͮT�x�I�N@�~덂t�_b��lw܍83�!�Nż�b��׾�0�4uP:���,b��_��io��_���h������2�u��dk�3�4�}\K��X��[��?equ�q��AfP�st�@u����c0��w�g=����+�Q�w
bsm;t�� S��=�ByW�AӲF�� �� ��=J�RrM���\>ڔ��daH=�8"?6��3j�J#6Y�D��`�@�t��Ü.�S{A�:�Ew�猶�����(��Y�0�g�����B]`������j?���x*�B�6��.�	f�� ̽Cjb~����F?��Wp��Mêe[P �L9vVͬ ��h&e�@�G$P�@?;�v���M�f��fI��#���bǛ��"���Y�>��:�0��Y1f�!L�:�JD�������7�nTx����X���o%���添A=q����ɚ��i	��Sito�Gȷ/2n'nZ��\�PEEy����H�k֑!Ծ� ,Ϛ ��:pĺ],U²�VsG"v��]U�Ld���&ձ��!������A*���Ѯ�V�A����dvU��_�0��u\�-Ch.h%��E���M�s��-�!�F��K�x*̐KjL��;�� ��$U�i�V�0�ai��q���2z韊,��P�%2ڭ9�����B
y������K)��H~*�FRs`�;:ٴ���n��LH$:1�|���c$8��=*?�1J)v8v	�2����<z�~&!:0ݘ��O˕3vrZt����0ȼ��:v�NUF�]��o��0L��JQ����Q5��+�����<��O��եr{m��&e��}���r����W1��+pT*����m���T��ϡ��١�J�p;����Ÿ�g�}�95��F�V'6�q'��͌�J`�4�*��}!�7�aY�H*kU��F۲%�n�#��m�6y��o��S��w��<c�[k�a���ʂ��k��a��v ��	�	C�"�����}ՒPˋ���/Kn���O�G�_*m���%��d>4jRk@�:V�*Ȥ*2��R �X�fa�K����)����i���"�q;����� =)u���Dar��0�D���6��E����l]�TDc��+�Ӄ��H�[��q*�Y��:=����+���� Ц�h���Ȗ,����8�ɦi��\����e#�!g� ~�y�1�ր��b�N�'���iU�+>^>�:�}��(�.^�ʝ����� ��pQ��{6�f$ף���^9�Z�OӠU��$��j#6~� ����9���B1�ݚ���v���	���K# P�p��逌��A	�K�����!N�P4b����7S�R�AsV��soO��0uZ9�u�pN	p7#�Qʤ�)�l8hA��fHE�n�'h�:AM��q��a�D��􉁒6��vlK�Q\���������%���\���gdI���T��ȏZ?  �H3�!n���؏��!>QS�=鯘tjR<����L;��䧏!�`/��(b�Z�r9ꬆ%�9gزN���$E�0�����?�=(��ϝYd6<e��'Sn�/R�txU3Ё�p���W4z* �>T������B�a;�녝�kX`�߶G�h)�!���=#�� G�A������imT��i0�n��!�T߆�N{"Ȱ�l�Yë,��@��Q{�?��v��dhO�g����[L����Y�u� ��Z��~��Ϣɣ���D��r~�����N�����|��3tpKT5�>n�e_D��D��+���9����x�ɭ�p��gD��;�aG�tx�n0ye_���W� +�M��(H��M_P��Z�jF����8�����@"UG�@yM���1.L�i^'���H74|���i��0���R�t��'T�|���t�Vj�R�}��@����?���c��=�;`Y뺮YS�Q���Al(�]y54��)ˣ�U$�e�PY�иDۚ���t�8�x��l:���ѕ��Y����!;�<�p��FR�}U��N��e�ɇj�̴���pϙv,%U"��Bg�K�y$ʺ
�q=��	�D��ax�B���e�-�
n@Q�+ȋ0[����7F�|<B�����d�;�o}��9�g)�h��t���*~5�����6�#��+����OU�7�$|A�a�9�`�3���/ F`"�/m�߅��5�0��p6n�u���OCD�z?�����-�2�օ/�S�~ƎIW����D2崮z}�ﴰ�eʱ�~V24�A�C�{�8~�tR����$�������"j�~�E*%�9��w�-K���Hsy�'B1a��r�����?F�֢�D����h/�FeR�"�se�5טk-�嫎r�b�B�����tS�][R��yR��i��m+���?��%9bJ��f�r�T��u������~���r�:��:~�K�v�dR����h��˨�q ���i鳊˲����1%g���>
��<�Ow������Y}ىqp����}Ze�6�!Kum??!>�0>(oF��ڑ�BSߟ<I�6����%�=����+�r��8�d>�������(xr���%-�EC�e�X;̩ܬPH|�� ����EC�pU���|~�~��b#dW���@_���']��+x���<~n��lʡ��O�ن%E��� twF������cYx#r�[Q{��r��@�b�~����P��b�k(b��v:j47$�[�=�A�K&����Z�c5��&���[��ӵX2���{;�Fv���%r;������^����\ka��&9������O��Y�������=��H�2��r��M~7��C�U6�W��&	W]��1Fd#���tJ���v��r�T�V�1௦w�ơ��נ��~��P�W�3S���#,;�VF�qH��n/���0@ә���ښ��]`�p�y�z-�������FK��+p΃K'�=`>�e���~��P먩�`C�Ra�Wa�ج	@������!��%�t��XsI�\)ж��6D�I'q�^�,a�/���M�#4nS��\c��%��m�1!����ʅ���n܈�f	�eW�ˌq�z���'���2@(N�<)]LG����`nJU���:ř�\k���/3�g�[�c�.���-�b��H#_�y#*J���A��uƏ\����%c��7x��Q�8𴁂����NN�ȑHnk_#��d���� ����4b�zPv���φm�%������`��P��a|z��Y��]�L'����z��[��Ρ�=�s���ؖ�Q9�Ha_��է�T�̈^����Xd�|���HI��wr��$/�����r���✃�Ξ�ؽ�<�_&�w�FU��f��x��[�M�^e	͉��j�?�OHz���
������^��f]���۸��*VB���ޟ�nv�M����lMI;}3��9S�}��}S��k%0�7�КJ�x��&L�L�v����˿����[�K8'���s伾�N�KϺ��w�@�L�*cpo�}ln�����*o�t�Ȃ�l�Ā@'�����Qcno5m����l���h��S籦�$�y�?7���տ���&&���2�%@&0U�$��ή���bT
.�+'���lmrB�\ߴ1R����.*�~C����P�|@E���w�_j��Kf��bu3�Q�Ae��&����{G*l����0.��I���	��~�-�f4}�gJ�6V/!N_'.����j��E=�W���`v�.��S����T7{��7����.���^�VYL�|:c#?;\���E��g�\#���(������@h+'�ʮY�SY>�Sq�e	�ٞ�+�,�4"jM�����T?���j)��^���¨)qk�.L�~ ���!:�Ⲵ��$�_'�+�잷Hy���q��r��r^�-�7@�JԔw*W����K�_�~�H�Q�d| `��n ���ABB6�oÄ�eѶ7�t}I�+uM�.���-�`D�x�q�n1������M�;�� 7� � i>�܇y$�.'��3&#��O�S��a��N�R�+s��m@07���W����Ը	�5�ُ����v�pz_$�ł�fɪRf�@�0����kr�+���Pls3ݍI�G�O38�I�Ĉ��b\��Ԑ�YdoUyA���W���Y��;-v($.:���-// )ӳEԫO���{�}(,�<��V.�C~���j:F-��{$|:���Pf5�4�/�|_��f�9ބ��JU�-�b^�
��E���ҵ�f|]==��チ��h��MI`�����_�9�?�X��wT�B�%��us�M�t4Ip!*��$6���	�錾�mIʩ��A�H|1�
���=`� N!��#�U�Y�c�ך.	��W���J�B�N��,��.9��C5rx��N����?�uҲtKx�]�H6� �.�Y��o�LJ|x;��W7�%ӟ')5+t��h�Qr�N��'3��Wɣ������hMV{6������u]��a�P��JН���ȉ2��f�F{,;۶w��M9dGئ�]�#��|�Ȍ曬ģ�4'p�G^�P=�� �ŊX�Ʉ��D������V��ف��M����P0�V������V�r�n(��H�F�۸[;Ȣ�k�ͱ�l��\e	b�2&z�
*>	IO�E����ػ��G�Q�刕"�x��`������A�w]� P[Z�O��WxzC�	�~�;�#Qelج��T��>q�6�% �_�4V��W��� ����t�v�חJDjm�%
��Ǵ�D�B��[�/�����{�; /R���ti�(�(Å�+��~P�zЗ�/�R��(�A\�Ϝ�n$s�v�%��"���'9�pzx��\h־7�j���a1L�!
����!�YX�m;W��k��e~q��W娮;8��/�E�J? �f��NB"k����I0��nB��V5�=��h���^�f�|Z\_���C��)�,)v� ��s4���Z��d��L�$L��s��a�%q�?��d�6�������B� ��bݧL(����<n�<}�B�ڃ��2��!�Yg��􄹰�n��rM�1���5��}�h�����l����v^?+�wʸ!�㞯�tg��M��M�;]x%�SR�E�m��&f�� 1�E��Z�v
�'JC�x��&�,�N�]���M##ᙐ(�|ŒO��/&�Ώig>e>|���O3=��֕ｶ(�Q��<@h-����j����ssv�1+����d�������z��~��)7�H3�D��Zn�͉aOa��s9��<�H�]}4�_���4v��sɖ�c��HŞP�Z�a��Wl���\�x;(Km�ϝ/?�8+��͕��T��kN$�^�!T��({���L h���C�|������6I�_h@�m���o�iV�)�/�I�ӱe�Wj�N��0�j�ȉ.�/]ǁU`��q��D.R��'K�ʐY��Z-6�U�� �dSw���D%��\}�"Եh�B�`�.�mR�]��/���] �%\+Xϣ�3CE����K�OqA�p��>�Z؏���D*��L}w���an���V�]�a�J��Hb�پ�[9�U��Tq�$������d�]ˠ��R�fQo,
'�1y(<����­�[��/��Rr:a�`̏՜�f��uޅ�jg����L�g˨�J�� 'J�It��L3Vx��yA. ��6�Z�\�c�Z")@�,�E����n@k{�&��%M`$f��q\%a��©ڜ�����{�R���/�~��(F�m�]�����뵪��z���b�b�śM>�����]^z��q���ig�3�\�*Qش��hJ���kY��� G���,�#K�J�>�r3L+����je
�r�OMĎ����xh�`�"�U8=Z\Y��}2j{��� s^)�Td	G�֢L��SL\Cb��z��eN��]�'"3���٣�0�F�d�$Q��q�%�`��ͅL'2�G��}2����;В�!��ABl�� J.bs��@ ��H�JA\bl@�"�z���Vˌ�c%���K6�����P���@  ��a��֌��V����I�S����dm+�Ⱥ$�.D!���.uL%���l��A&V�6�1J D��U��P�Т�ܗ�b��̹6�����CD�i��,NMl[aB��n��Л�Qϝ�����G�!*��3��.l��8٬�r�P�l�9XE3��>l�ध}�A��7?p!�8�U_7+���+���T5�5�*(������[��zz2��[�e��m�p�����z%wMz;�z?�B���9b���D}G'oYoUȎ�1�����U����X�N�g��"(3_3e�A}h�Y�0�b��&3�C��TGd$��s��#���{!T@��|��L(7=sU
���=~w�
���?v��*9�#�X�0����(��9��پ\�)0$��샶^'�7�tR-��C�*+,16���di�'���z�Y�١?�V%DDS����l���(ӂq����3i��_Vf%�Z�8�1' b7(�. �����Z0S|�W���f/�d�B����U7��l�W��9�<��o��c�ʶ�E�7�1��²��Z
+�_�ɴ܋�>���[�Е�r1
�)���f�<����g&����C-��v��Q�b��X�n;�fۈ���$i����D�����ܴ�љ�j���@T-��,��0lO�' m����o��u@��o���oy���"#p��A�EA�\:�}�
�3��P������7��՞{c�(F���C~dh��M�S;��C��lh���֪f{I��E6�����:'0P��F��d=~b	E���:�R2���)�6�\�
�U(}��b��ك@(�2�����%پ�������l�T<���:��ˎ�P��/��q!�o��r���F��HŴu�ǂ�jh0�R*��=�V������[`^L>
B��Ǽ��`X��p�_G��Xd��Q�s�Q+ly+h4^�:��tӾ��LrI�S�->y��ܾ"�o����5�����w��N��O�B�������G�/�m�j���Ѱwc�Ram�oA��d�r�KvR�bRv'�.�k��I=�j���ܰ�`*��	�Ĵ��`1_��Ɍ�����R��݊��C���� ������m��FE��!��R!)��-���ݙE����fL�ab��#+r�[����h\����䍝�w�����ZS��F+'���k1 �G�FI��MM��#��1�d���a8��<���C�57)i��T�q�Y 6�^MWW'����5�Q��%U<F��ї�*��	=l������}�\;�s�R�!�ѵ	������S���q�w�P�i^�UXp<�e�hކ�,��P۟�j~�%?��#V��v��G'�FMYu_T.���6��5$"�9�bw���"�Lyp�T�zT��%��{7�9��� ȇ����ý�4n��߶�2'�
����S�U��>�oM�hR�.|�9��,�E�����mq���6�WK$L�1��*�0E������hd� jk�Y�8;��:��h��Ѩ��/�D��opˢ.ɥ/��l(�_"l/$��0
wx�o�'���(���.o��"y�A	d�����"�����Q�N6�m��2����6,�������ޔ���[e����.�	Q" =� ?#�c�dtY9�H�9��Aذ-E��x��F�����{s����K���9Δ|��@~O���e|}�-�X�Q��|(U��=�"�Hr��'��
�Ng+��V\�Yd��7��02�~_��Ӌ>��?4-��r�?^�	��w�ߖ�È=;�Kb�n��I.A)P'������>x�A���7����'Nv�����R��=F�U���� ���f��A}U\l��)���lĈ/��!T��~����.|�Z��)�ØV-gq�
S�_3?�9�|��g^>��/�h���B��7�}�}�3xl[���[�b"Yy@�T����$�;���(�$ֻ�I�_�.�T������B|[���˜�A�,G 90Gx�2��+4�Q�Kڍ��=��qŽ�f�u��+���B��B�nMJ)Tl�;Ř39v������7�ݹ}���?!�����p�D����ߒ$S�w�\�LSC�Z�ov���]��V�G+�F�a���.�Q^�/����-W���֧I�d�F���:m���8�j�Hl@#��Me��.ؚ$ax��{��6#��n���g�e�+���ix���+d*�����뢕��':��v�jO��D�BF�l��x6����eR}ª�rb���Ǩ/9���j�*�:i�I-��}��op������_����Ql���*r�@r�CdP4B^ґDQo���qm��������_�a�@6�颚�f�A�R�B���is�U�=]��2���O.�2D�>(`���	�~�� ӱ����m��xif�P>F̠a�M�֡��nq��6�j������WQG���B}]Ǥ�QA��?ۂ�ȸ�EV��x>uʘK�Jv����F�>�|D�+�z�x
E�/��]wpkH�JUX�%�3ȥꖃ��* ��(��C�<4�e�5*����e3��?��M"#3MgM��{g�g������u4��4�� �㷐�Vd�u�m6�k���@,�:Fk[Җ7bQI ���s6]��{���I�F]CT@��[�������-R"�l]�.���!�4D��BR���`�R��-%����ȃ~�4'q���s��O��Aa�h臃��gX�n��$�OΛ����s(���ED��"�#?�,�Z,xRD��+�G
#Œ�"�0u���L����_t�+�c�:zM.��D�֏�ۛ��k�>��f�&@���37*IH�^+ܮ}��T	�^�-�4�a����S�Yi���ɱ:��8�W}`׽I���Yr��<-쒸��Br��c[���^��>�Ks�c8oҠ�\&��4R����ߍ��8&7�?Τ�:{��Sw�V��	H�ب�C�9�9�'�
��T���	o\՜l�kӇUe��ï_|&�f�ݑѪD�*34ݢ�hҮ���A����#��3�v#��B��;�1�Yh��#hnGFցOKP}�A��hl����?�=��է�l�!�I�'q묎
^�� ���� }��Ի6˙��-�M[�8�\�hB@�v:�y���K�A���[s:~�<�%����|o.�ᢢ6��t��q�xg 	�����p�"R�+�@Z��}Δ�&���u��,����݌VM�#�(�����CI���Qqк����+���"b������o�&3L�$'�Uw���b� �w`�0��R {a!rJ`������f��ImXwI�z�f#M��a��N�wA�=�R����l��gO?�] �f�ٽ�jǭ*f��+�sҐ5�������_�񎱃�+I,ԙ�Lt���'J%��q7��c�謊���N뉦�
�3����y����T[n^�FHN�)Ӱ��s������!�rg�k7�呗�z��i���H�k���~_]*��~���s�O_�Li�4�;]:HY�",?G���	>ȕ�ޮC�����G�Qg�e�E+�U���`�0�@���e0��w��M��:i�^FF�d�(j�st���n:_w���
1=�1��	��	L��A�"��e�6Z�>ja�_�J��4p6Hl�YF�܄��"m��; S��f����ؐ&���QYeD �ˆ,�P��rY��i� 9"��B�}J��?x��kZ+��d�-]�	t��0z颲
�p��M�jpz{F���3⹅����>ڻh;�a�zUT�T�)�$(w��S���
��"�]v�q��֤?���)Nn���y�*R����m�e�~���<h���X�e� <C�obz�d��ݚ��z̧ٴ���Ԍ��s��#UX3�f��/HhK���+.b@�&E�
Ο:�U9�:�rU<[�hQ�m�1��I��f����>r�<G�����hi�*;�e�)�7��-����3;.����	ةiWpY�C�Aq�!��M��?��x,�h��ڕ���#��+��a�=�[	� �JҮ��q�ԅ}����,�.��ɬ;#�؀���W���R~1W���D� ��i��FK
q�(��L��n͛���|Ή[�g�w�0�7X�l��z�h<Y�K_��B�U_6���V��������ztN��͈~�nB��fBͼz�+:#�:�ܔ
���c���i���!gUGg��s0�C��1:�N�5�M.?:���١��F��*$|��y���/�H�qP�����@2)��VI�26X:�{�G *[J�`�� � �</P����;o�-0hv}�2��\�+?;�ϋ�r��-���k�G�	/7:�X�I-4���8�2m��&9��I3CKQq_w��jQRӮ2���a�rӃ���+#ޏ B�Z�MH��'�:.�����3�D�
;O"\q\Q
��te����	1ЇG(�{�!Xx_y.6� I�^Z�iJ���5�%���v��g�_yrG3��		����S�`���	4u�Ʌ��׀z:�V�����%5�pc~<FK��íBΕ3��<���Մ��@
���}���\{��x�c�-�����Eu��(m͝$�c�]�����ވDO̗�'�1�7�l8f�T:��_��)GV~�v�-�e�7OAp���(�W�~'cf�U��	ML�)H^f'��p%;mp^Ӛ���z�g#�����H���b<�����^�?�θ�A��/�F�R&=f�n��l��sc���i��)�9d��d2#�Y` �y��X���^O1M~p1���b��R���/����u�Mo����J�����>��o���Fu�ΰVEeR�T�����g�i�#�xM��T�fƥ�S��i�gadA'�l7�l޶ �j!G+]�iZ��`yW6w/&P}Je������^�s�vG;w�^�t�v��dѐ�o�8ug�!����K�ɔ�F���0��}[K5W�j@E��?)_i�͞�|����d-�0-��UݺBgb����yw�"l�����ȧTZe�zPC>u\��Y�Op}�;���M2��� 2�X�9z�� H$bPdIc��:� n3�)*q}�,�i�p���덷!]~��#���x=|�|I%2�K�~iA^:܇c�SW#fj���i�1���1~Mo�-^�02�D�]�.O̢�:����MmT[t%�`��y+�|;b]ב����u��ƈn�y�s��tMV�"��|�̃l���>�6�W�;�R�O��jpk�|z{B��<���8��:��
��mK<����_J�<�>�E�4[�׽
�0(�-v���sWt;;ό}����^\��ox'=�w�5��-��%J�D���#�߼�X+e�{�"|���q
����M��H@qWēk�K���n^��:��z�X�_���%���.m��x�A%;#D^+{&�՟�ͨxχ,ӎ���I�C�!8��H���q��8�$:5,d�x��������Z�z���"�(	���$Tm��:�W��-���KkP|~�p�l�K� ���;���=f��o��V&�k�w��׊���7����M������:/���ӋL�v��S+��~��c��R`8���v�	�8��{~.˧�dN�(�8^��q��R�~���TP�y2,���o�(u���|��p�Oc�h��i����y����f&�#nKH�_�¸�3���눡�Y�u�7U�����Y.А�du�MSYv�2z]�)��P�O��qiC�xT7a��K'kxGt��BW%���#G���>я��O��2!nix�Ji��߯hG�sgg��?j=���d�S�[�hk:I�ﺃ;��3Z���l�Ĺ�fj��h8J�{�(\�>N��y��%������$=��E�͚�ɚ��=��-q��6E�
�ՓN�@B�@i�8Y-�)(��Så�B��1'��$i�O�g��Ӻ�'Ϗ�a+4�fAr������+;�S�����w����c�u� ��c���ZX&�ߍǬ�ʔ�ͭ�&Av��{�g�a��E��1ql(��Or?iK�nw�~n[7�^C\|^�����ɠ�Ѭ��jf�a��u��f�P��;��_�D���%Z8l-Oe��!�>�0M�p˟�8g�5�6}���Q�����@-��]�-z}z
 k#GTd:\kˢC��Z}�0��O��_y)]t ��B;:�Ս< �m�(������u��f6�A��.n�f
VA� �'҇g�����y���iw�����b9�\T���_�
����/�P�G���;��9z_��8�?�46��0�E%'�ϫGd�!Z?�i��}s�����ln��g�*ж9x�3��x؛����T���On�!G���r����Pֳ�(��Q�e⺺���c�j�u�N�r��i��=��!{���z��@1�Egݭ�fܔ!Nﭓ�t�y <e$.r�S��s��?����K�h��3�n���4w�'Y���;�|��vU��Uf�[���@!'z�в�S� ��nӆK�}��Ds�Y=?=�%���m���.����Q�r�9�&[K�G�n�����z�oL�걈Ɓ��{֌�q�ŗ&/D�$"�V�F�L͂��י\�"�c��q��E%RJ�WA}AY)�����qH:��a��)g������r��ss�aN���)�� �ϻ��/Q�_�n��
�?�ȋq�I�
ӻ�s떣�ɴ|�8D�I�z��|yN����oI�' �N�-�;��T���ZF�A��[�����ne���>�&�s�eѵ����BZ�b�����;n��-zV(^�䆹�A�b�N��M'����-��S�*jԶ�ݡdI���@է�v��9��d.:����PHI��_0�-����,���?��<4 ����H���Bi;��褩�(�^�)��J�`n`�[Y&�ɲ��eO+]��ZW�)��]@g�IC<Yt
�9s#��2���H�_xZH��e���*G�l�C}�Y׋K3���ʟɉM�}�=݅r�m��Ψ�4����wR-襠���؆4�h�\Δ�q̔.�q�=4�>N�h��(��T8�]�K�P�d���.�Ͱ=o��՘��y>W��x0*?��	���Bl��e�<I���w��`�B�g �`�/�����O����W���E�����=��绛�-#+��m��AtMS��H�V$�v�
G����oݣ����w�g���ό�z�����b���qnNf�*�ͽ���E�,��m��	
%kRH5�s`$18�0�+��uJѼH�H:�<F�� 9�ϥ����#tDؚ�����ȥ��Y��T��Hl�l�¸J�G�Z-Ys6 ��^����l5CA�"sVBR:	���Ш�#�r�Y1�ʳ>�� ��r��m���0c-&o�[_y�����@��*ѣi���$�%�lj(*�K;eҳ�Q6g� ��9m78'��OvIrRB�~$���G[���~Z�|�[-�{CnS����]���sO5�<��!�A/#�����'�Q0t,\���nw0�^�kSA{o���sF|��)
b)SQ�'m&�ψͪX2R�pkc���A��z�c�����xū�~�{F�����8�hbw�]��3��-?�������x훳w���x_`�i&��Ə��?�S�hPU�ϊ��^v�ś&�@8�R�n �L#�0PE��,��9��YИS9��9fAg�ᡂ�Gq�.�ႿP���<`���#7
��*w����"��Vl3/����[��t}Qv�D���pF0N>Q[V�Ȳ>AG�c���k|@?@Z��ãg{�{��)�\V4����vYY�ǖ�����(p�־1]}��l�w�X�yo�7ɦ,�o�/����h��)a�2�ܪ7��`�"���%�����ڃ�N*���$N+ )q�m�}�M5څ�h�k?���<�D�@5�u���iY��K�1��E�t���E�wÀ�x��� Β6p���
Q��*��$Y�+�h&Dqr�Q�ow�Q���t%;�|+]5&��c�SYN��مVaR�T�Q��(���V4�2��^�_�p�7ɥ�+,�ך�|QK��I���i�+z
R����|�����Vp�z ��}�I ܏��$G� ���"G�sſD�=5-�N��O�k������>(.��֨�'�n��-��
Mb�JX����0+V��ka�	>�z�Jigo5�����6
���z��� ������2��ZT��1��������M��~�dS�E��#\���)��P|�{v���}C5�<�
���ݓ� V;5�FR�@3=����d+O����C�ʳ|�AP`����+#�5W5ݗ���0� �S��T]�:"����Uy�����< ���K�Y�=�L����[z�)F5��v�!/uL4b����hMlw�U!1��U��;�x�{�i����@�9�>v�����N�[���'�G�T��R�C��|@�T6�����a
�B�G�zF�Ll6EW�|�ʧ��ա?Lfg�~��i�e��P�~���7M���W�O��a����NA(�%D���������&�����@�{ @�._���������ڠ��v�4^��	_kYTD�&i?{��8*���9;�f��|�f�w���EvA��D(4W��H:a���A䛿a�P�傠�3���J��={��J���(�Y���KL9=��0�<�� ��pG��.��qUY0E�d��6��2=�)
<[�@L��R#4��TX��|�Yϛll���c(�= � �\��*�7y_��~r��w��	(n��ԋy���T}�I����Þ�i���{s��)� �]I�θ�M�}g0�~x������Tq��+k�'��
�M�=�C��H�5Z"R�+.-��(<�矁���Q�E�$]$l}�k��@]��k�ϱ��>|J��8���ŃR��c���E�@����ҳ:���
���ի	h�8��O!��iO6�p��DIw&++�$w�Ѹ(�;�6)'n�VHt[�vj[��i1�x�Z蝐���P�}�2>*�[��X�ݮuH<�c�b�L	j�	�༝}���B���*P�HX����?m|7B�s���pwv�W��Q��I�)w�$U�E���y�j"&����^ ��v��'Iʟ5ݷ�z`�L�����s�K g�5]^�J�6c�v��"~��(*Q�� i���'�����[A��"�8�D+�߇�`��_J�Bl��7B("��%'������]2���h����/ �,�?�z|���2TF�3$�g2�xfu��k���`f0�]�Aa��6�-�L��n��*H#Ã�o���a-n�B)�N��Z!xc�?�\a��_8��ڕ}�l��)
�,���6�'��r=��멸�����4M׷SU���"r" �S��$紱$s]�`��/-yʹ̟1��<~Ym,� K���
r�+&�������S���Cg�r���-�=57���S�ǣ^mĠ���|��"P���UA�=y��Cɸ��,m��� �����< JY a��2ܝ�
o<�R1=X��#*�:|��� ���j�	IR�N����+��/A!|Ո�V�^Y8��J�V�<�$��_��X �e��g?u���x�J&��hq�'n�@k'$)?RF�`흤}�$�jw�����9u�[j�NgZV<��o:ʷ�!~�# Ezdhx�ܛ�'�����'�����H��1��ى��S>FjI�����Rc3��_D�Ķ�͖]#���3�;�䀹t�T�_�������Z%���K��h�.�E��q�j@�����е�� {|J��MkaO���&�U�A�n�w��k�:��c܀�{�W����աh���D�UGR� N4��24k�Է�|��o�<�0g����=��gh:Bk���Z�M�8'w�C��`W�O���Jl=��m>`�����'�ԷseK�����i���h:��|wꃟߘQ�9�B�;2곿&h�p��(�ML4�#�Y�O[Z�J�m7������"y�[)@�l�O[-˘g��h�0�0(Q����ǹ�<߆4E���|��q:9ȚS��w��}Xr�Ӳ�ܥ�I��av�vȓ1a�[̛�X�H����`;}(�Y�͢lT�.�hY�-���P�q���;�9#m���H8'6m,� �N �1�W.�K����,�����E��)yg` }+�過��,�}k�!���@�+�����^ 淲��������i��'��h��Ꮋ�{)UN���w�5�!��h���6�)�4�b5ۘ����ɯ�!	��R�/��Z�Ѧ�d({w?�Q0�	��Dy g7���g�Bu�)O�Qk��$LZ.kU������_��;�8Ky���x�S�!t�>�P�3�NF����Ή Tx�0Bwq����
՗�!��m��.��4c�=�餰����o���l0O��g��w�;`��|�UPy�ε<�RO���@�x��kP����Q�(�^pu{�����gh����d~x�f*fv�똈"�����A��q9�7!�h�b)�?dd�Eu�X�B�w�d{��Z�:�\���g�!��y�q!�k���~#-X<="z�JU��A���,��'�;����Z�0W�w��O�F�k����"K�\5H�#�:{�xu�D��F��1 y6xC-�'3�Zy��H:"B�{	�����ZA�f&:�6'��?ބ���V��ގ����ц[���k��0�6Se@�"n��9����)�w����;l>�Sb|ԏ�Q�r�(n�b�Y�-5�0�|S��L�0�wAF���af%X$]�f����Rm�m��!�'�\a��Aş�2�łNc���w�����M`˦�ԍ���4X�S=bK�F�Y�je	�$)��B;._��(���e��J�j�6	��SC����^ϑOՌ}L��-=�Ӻ��Pu*8n��tka�v��(���[x���>�� =$9�)��p���,%��[ó��
���M�:7�H�m��Muu�]`]�Qw&�mG&���'��� �����j�{(��t�JC�Ÿ���I�<R>�5�`좚�I�B3Dc֨�u�گ"�A�6@л����(+�ö�]^H�1d��=�OCQ�}Vf�����/��'L��x=2j��Ӑ�����r"8'�.����B ID������N��r�݆3���O�ʧ��mv7;f�&�I��ĹX�3��G��}��REe �KGMap�d���5l�X��П]!���ݲ���Q3��O��p�Yv����8
Y��dlsog�'α+�)S��"�H D'�a1P�5+:��r`�I;E���EkKg�I�(.��h�q^��d����}i��m�δ��K�p !�W�.b�r�	%M��Vv���.J����^�t���A���-_����0����.-��,��K����D���8c�6��K��l/^v���4yvnV9�S�����s��)��N �y5�__��=�i�"���5cۼ�Q����`��|�Y\����~s�;an[�|Wz=	!PS�~ <��{�To������CFd)���S��-'��=5��w{C���w��Ы��s>�2�
�Dݽ[�!��^Q;��WR�T��݉Z�_E\��Z�D$[�N��4�z�#��_g��a��F����r�����:��A�_��Z�,=m�$yf���s� ����ya�s����u4������L��D��ο�7P65�a���$�:���QW��1�	�Gt{6���2ʴ//�d��aqjqn���+�4��h�Ʈ͆�ߖ(Jɪ܇Q'��2cEm�7��4���X��7T�O
��>��Y����Z	���\����=a_�&��|I�����(��I���E'��\�E�W�#�ci &u�T�;���=���A!��%��W ����Q��횂��g�:0�6�o3�-v�/ą��Cޘ,�Pk�y����	�����.�,3� �~�N�����@�s2�5l.9Y�BIu����{�yG������Q��!�U�[�_�������O�������@O��!�<ȭdF>Y0�5IF��C�&��M��&�]�k[q���찀��V"%u�5�̝��?Ca��qU��C��Ys����<w�4~2��	i��R��La��Q�We�E�U��X��_hCu~�]���7��ӫ�]|Z}F���)��5t^�?��=��F�b}�*#�i��y�1{��I*R��l���"�1(� կa����s@��e��R����VQ)�~��x�ޅ�UՁL�9?��N�iM�����ޜwb�
�8RqcvIoCy�hu����ː�`?�(/�W����������k�e���	��!�yX��*!���>��S��#"�CC�X�������v�4O�Me S>Jt���\�Y�¦��I���wC��`���[�����o�v虬�/��V����|�=��aye���iوܛJK�qP�(�x�� ��l����v��2�SZ�t <�G,{�,�7�Ⱥ9���p:*�Z�2
^L�»�>�����=�"�m��e�]wӞ�y��LN��N5��	��S��I��*�/�m�k�������2=*��"�c{��o��~��WˆU��|*o��Zp��.�I��Yv"T��|��tb:�H8�Q�E�
��yϸK��~d���cs��e�s�_ \sٙ��f�i,4"�YٞWaҺ+u�+?َ���s�I�m�^|h�I���
��P.Y|���Z�h��~� ��x�7]�J�x���y�m`M#��{�5h% ����b"(���?��x�K��C�-/{���؛tV��A7��ŭF+�0noX��k�=�8�Gϒ���}/?�f��!.`t�C ���N%�R��4z�@[��)�x�+ ���!6��^�i)��YW��P�'h���c�@8����S�pj=��\(�c(62��2"1�>t���`�������{�L#�`��^e!R�2�4D��n��Fq�v�V�m�qX�Pf���KG�R�M<�~�}���7�����?��N��ж�8������!B���t}�L�8�.� 7�e�FEq�����V��\=NI�y�-�s�
Ƅ��z��p[J��8�b0q��W�Bل�R���Obu�r�f����*���2�%̪<�0i��p
�3
G�8����Q�r�k�h��f�$Z��u"ɞ��:��y��ޢ��HNn+�� �6⬵͵��^��X�e_)�jb�>㒰�.��X��j{u|�%j��i,U��Mb>��a:����1+�ګ� �W�*OCy����u������~�e�x<��1y��MwEI ��Z� [g�[;����M��6nfv>c��LBH���8��p����N�s�aWZp�L�XO�U1�:���J��띗����?h���(�
{�&�[Σ�?o��|?k5�?�d��Ū\/���H<s�$��+�p��ǼEB�7ʮ������X)��H�-p��P��ɎRcf�_N&�u���[�d!�ٜ��ȓ�[�}S/�o8��
��A��nTjyu��N��־��0������T��G��C=�z#��|u`r��W@�J�V�'*���ʝ�ъ�m�����\*��f��$���_��+��Ie��'���ƾbQ�q���=b_rͶ;XB`&i\��GX���jR�����:(Εʢ6����a�����S�X��vXC̂�U	�V�E�j�����m��u�`a���0�E�{��g\�T�a��{ɝv��\;F{�3z�/Y5�ޛ0���g��0�Q��f�؛�6<A&]Ś�,�q[�!�ab�-�E����}4�kuaߖ��pz���SV����07�`�������z�t�5G��;K:j�Q�[5c�Em�D0M��^�aYܪ���g�^D�v` )#�!�ms1K"��}]٭Z-�|�*5�At[l�(k�˜m��_�R�!L��GV��}�<E$D>5#�u���hK���'���
x+�p%q�<`��a5	i~�!�r��7�~��A��c�Q}��QSd�s�7� �M����>�� ����	��gR���X��8qE�ӿ?�*����xY��[�>�a'ֻ]�z�DGBC�F�\{�Nx�qr:�P�龤��H�d�/P/�l�;ggs�MM

a�-� 2o�( �HP l���N���f�+�O���H��)���ؤUl��d���(�˩���A��P�fdl���v�X�q�Q#w3M�"mrU����%s�oei>p��l���/~v�ǿAH-�=��U�O��L���J8��*j@�|>��$���{�)�Ak)ܓ�6P���v��B`���R(w!��4��v�?��9�+$�b��w|4�Fp0���	�%�	���`t'*�P�[~��Kag`��b�C���x.^튣�K��9љ�'�ߥ� �'�0.�s3=IO{*w�t�~7�ְ�U����޷Q@0_��Z4r�6u�B��p��2����v��1��P#��s�@�����ؠ0�_$����(.�c��S�w_F(t�6s?Z���ʪ�� �UQ0��Z�$N���`4��E��H�nSTb'��D�/*3�7�{��p���got�t� ܣ�\�hO��f�q� ���c�t�2K>��T
��m����4T�X����l�~T�_U
 B�!��Z`X͘���)�8YI���#@��(rG�.�:�������(�(�5��}&:l��S�b�'�,�_���pr�N���'���soE�7�fM��4L������}�^ 1��H*�'=��C�Q��/`��+��b :��px��ܣzD�B
c���K
����]���s���u��3�˽}�*$'�� �>��cm�����Ĩ�S4	���˛<`E���^���^:�Q\�6����E����_D7$���@c�w2+M�D��p����:�Oz�Y�Άs|�\�>Ay/�8��@u�&�9m��}�|�S�36¡�dH�:`���s)Q#ؒ�odBx��S����8
��ȥ	6�0���@��F
f�/!â�����b���5o-�P8^=�q�)��:4�q��Y/�_�b.�M�x��Z;ǭ��m�a"M��� r���9|���ӄ�"���%3,�k1��,7��9�)AgX�JDka%��H�ܟ�e���ƫNU���9i����r�m�=�<a����іQ� ���ʝr}a�[��ɕ�j�* ZL���:�����`j��7B�g��2������<� �~��/� ��b}�:)�/��Z�X�}��A
\'�:�?���Xr���p�U�/�k}��eZ�|~��e#l�Y�q5�*к�s���u'��u��'��D��a�JDIO�c�bq)����-�!,�bm�ui��	�*Y�F�f3�x�*3����%��Z��}9��/��b����� H��Ğ+�>����2ɑ��ҿ�Z��49"�m��|
����t�﮸/���g��
�7:���κ�˩cJ���7*��%�$[�c��e�����&|5���s�k����9CE��8���7�,�	p2�����fE�zC�p��o���]U/�L�k��ѲȵL*�Q$�;x�"�0��կ�1bYX��$V]����B�	�ř$b�9Z(��Y��
%zh�RS�2.���`e����o�o� V��ӝ�����P�x�
�	q	�9�"x'9z5�p��-���S��B���I �Q:��	#�������e)�R�_��k-E7�ur���/>#6c ��6 �}�%����m����h;�5*?<��7������_"�}�88��	����@��MK�K��w��lW���l�=�ߎ��J+���4��?�����HJ�D5
���?���K�5���8�4۪tU�f��V;�,���<���7�D��1��a�-��Lb�w�|������Va �.��f��� �B���ȪT�A��g͑��'�$D��-_��;[�8ҶG�$-�����+�丌$��_�<ɴ�7���N��O�3I�.�TҔ܀Ss��v�cL|ZAj�������Y@jj6٘���Um��tsN�8�ǫ^���3j�_��R=���{.�qb������Ρm�B ��ޛк����� ��B	h簴��zd��=�C�8�Lm3ݬO1�-��o�U�J��ς/�?�C�� �/ʫS�ݪ��뷩S�����tD�Ώȟ ��y/��C]��r�L�R��׾pc�~�[ü����C�Y� ٠bY��g�t�U��'��F�,��ӂh�cM������kf�pJ$�ŋ���
��`�A�H��P �l�F�NtV�4*j_�UZ�\`��!�8*�rS�N��q�P�)\.4bԱ�B�\��:�L�%-SG@�s��4��Ϧv�gt�;�����쏟K��؏�88f�n���B孕��cð}�G�5��%���3T�ch}����� �,V����)a���!NV���X�eb�!����_�pu5��MȔ%�}aq�_�Ӳ��q��Y ���ɥ��]�)�b���$gs��p�cL"���-�1�G�J� ���f)Ҵ[�q-�'�U���o]��b+�9qq��Z��2���^�#q��-\���hՍ�(f����&C�v��`�w`QI�i�Veظ&��7��$~�m��H�b���T�s�o����������7,UgŰ�`�����M�����1����t��Qt��vxa^���k�c�]��/��w�1�I��6�����si;N�H�ofAW�O�׃�14���WH�N�������!���ˊE�ܩ~�͢�B�����r.hT��Y���H�a�=���]?d���]Q�%%-��]�]3��Ț>�~?�\XG�s�`�Yoqz�@�>�n+]"1G$n�7�+�,j�c|ƞ��k|<FZ�{�L��Vb�Hc�:�*��=�����Ʌ�n��qp�5ϧ��@.�:MO\�{��$��J�o�����.)2eG2��`*��� �0�*]:~��z�7�&�(	
�e�<
�K9Ƿ�8���AsFyA>����|��` y�FRyW���N9�M�ʏ}c	��C7l�S
~A���Hc�j���{}*����$�=+l��YУ�t\Dg��{p:��O9<��\<�v���������>�]��i����z:�թ}@�bS:'���޷ץ�����{�mcq� ��ׅ�x\�%��W,���_}���~�qZ��S���!��)�"����&3t��X<\�o�V�J#��K�`_܈�$��z���٤��q�G�19�d��qᣆ_F�I�h�g�<m�7o
ʛw|��P�/�J�P��z�Ӂ�a���ü3�@�? D��fyg��	�=�� uW�ç`�U�>i��S�J��PX�p�x@Oҩg�� ��c�kŐ��u_:�ѷ�["{��챞 ����W���l:r�����C,��į�*��$����4{2D<p�����Gr�2�~Wq,�;������������O(�>)�H��s��P�ɳ�R�[-5fB*y�
����n�T	b�p��=����<]j[>&!��^�O�>o�L�,6S'D'��n����o�F+����e9GO�� $���v�ό�1�w�����v#f�:/R�83.�v<��w�۟�.�OG�*���/���7a�,�\Z�_�9Q�On����ɦ,�}�����2j8����A�kk�J�9��
T�ێb��AZ]'R�O�:�B�nmK�}J��{�v�(m<Ȣ������]f�՛��o�y���!�p����%��ކ_cR����,dh���m���M�6�G�o~�����\B��~7u/��y���z*o���ʄM���g�I�+�:χC�-n|# 3gڂ��v���>=����3 gY���/:��`���[��y0��-6���*qjR,E�C�> ��H������q�a�>ǩG"j_�2f�?�i�F.�njS$UI��+��>�.�M�N����N�H�c\�@ �N���Y�2sOL��C�QUI؋�}d(n*�Ht.*��;�֌<�w�=8fb��',&������Qb^��':�����9�g)�8�ӣ_ɞ|���;猼n���c�d������Б����p�g���u�<��/C��tD���Jy��Q�~���L������5g���zSS�� �E��k%��i�|X{T�3]o�*TD���]R���I�N�>�D8J�����ЏT8klQ�z�#0�đms�Y�aȮ� w������o�ro�� �K@�5XDé GSe�&fyx�d��
獚-������������x���=�<c����SJʚV���L>�3�
����4���H>cl����l�k1��־�|9�������-� o<��8*��y��QQ�3�0��|K���c
�'\��bq�&�E��tX�6���G/C��1ez�zETT�w����S�g�+:�܍���z��8k(Kw�,`�1�*Q�2 �~��[Ɍs����B�n�eO2S�������_�� "�o4`���<�q*�XV@�Ȫ��1d�9Q�OnMKL�~�j��LT�&��[��-2Bi�Z@��f)O$\�doX�ZwP�A����ī�[/�����"B&p+՗L �g�e�' �b��Vt��;��J%�)�;X&��9l�`�����R 6}�R�"�V���!j��Π��l��� �{�:����HԼ	?s}Ed
3��S�Dj��׬yA\&��짝���^�,�׋�1���f���6WBf0�//�UOv��H4{W8Ľ�S�%(��Ģ�X��tC^g=��ORj�VB�����v~���"�ڼ�!Bt]O,+e{�$�F(7U�5r^�~��,%�
��fdk�&?�*�`���oQ���*.\�Nn�OJ���ǒ�T1X�h][�X�,	J|UiwL��E��\�3�����ѡcM�Oк?��:�T�
@�_1��oB�	MȤ�s�h��H����GH��·����\FrU���㺋�x֞\���)�ɇ\�s�S�[j�b��D#�H-��޷'3�b��[�<^;�1ӿ%�	�u�4;9�Iƥ��i�����HĹV���E��;�Y���fU�ZN�O�3�@^�ٜ��!� ��}�*�u�f�Y?���u�.lJ
x�6�z����}��
0_��ТI����)nx�']XR3}*�%�?�����[�i�Yg2۹Qq���T��l��6o5�;�D��x��wZ�u7����u����[?�7:�m�f~Y`�6�,?�b��ϵ"�*�&'�2�e��g�5F�'y�P���}��^��M<���o�xr{�2d��ɍ^3�`S/����7�a�G\C�G7sp�A�i"��	%���qū�	MR�ຎ��9
�8X *OY-.�KF�&��<d��\��	����J�s��FN���_���'�9�a�p�=g�5vH1��=!o�K%݅�N�����̤���ET1Ls�6�?u�Q� <��F�Cⴤ��F�����a���П��kE�(61Kٷ��[�\���_74ܥ\�H�9���9p��Y��R�(�>OcuO������͂�y�/3��⯃q�n/o.�L��q�b����O���{��r�g���Ä�?��s���*��h)Uז�]���Ѣ�y���`����]��;w(&�[ǒ��8�P*ѧ`�1Y�P�w�,F_&�<��;�������.s'������FeG���,_��{Sݎ�_K}.e�:5��#f���F�Z|t�x���Ƹ�A��Ģ��|�SF*��'r�i?�i֨���>�Yk���$?GcX�NC�אt�Q�t%�-Z���c��e��B�"�=��1�㮈�D�.�����.�_���h���I�df��>�c��/۰
k���{�D��è�����XG�m�mP��)�9�.��æ�c���-�����Jʓ�vn;@�P(i�����3	~�٢�/TPs��j��b*F/-	�!C��Tg�A=��Q�vC�<�������s�D3�͋ZH{���E������ʊ*o;b{�:��2=����a���[?�t�J>Zժ�f!�O�uH���Ofʆ+���J0�u��Y̻�c��i��z_�Vр/iWxVm�KQ���>�Il=�~��ؚ	-ݽ���+���������)C�߆���q�E����	�@����p^T��u�G>|�^��~�/ J)��nd�t� nQ[;7��Z�عǁL��z�%��󫖃vnR|
������%��j��ۺ��*�:�e�v��%�
g�'vV6��]1�@%o��O^�\���p����G{(�i�4�br���)�^س�?:�F:,��&Pٚ^X�)_ث����a�W�j�`qm�N�:唽���fr&�*�i%���_yFpp���E�V�;�	h&���4��YQ��?��$ܹ�u�
�)�2W7���j^��q�bB7O����3J��b�fq4�C�%c�o9�x�J�~�|}�Nu";+�7_Kp|)xJ&۾�O�xxl�3)E�����)��ۨ�!~�7�[�&��gV�͆��%��A��];��i%=AP�au�U��nS���ԴT+X�B�ҭiuM^����]��J�?��ޭJw[�M�Y��o����7���GZK�k��-ΌfĈw�`_���W-�7�e"���Ǣ_��"�9���_�,�h�'��u��q4���8Flf��]a���;0#e�+՘��nh�����[uSH�D��c��v�ݡ�4ڭ�+s&�(�q�a���塑B�2�b��yw�ZUJ�'.Q��h��� �����z�;Y�
�`cuP���GzԼ	Y<╧��
4� �|6����YV�P<M|�*��ݶ�<���/�GgMu� �����\���(�R]O����$Z��snņ�zo
D�U�[ ��X'�;�lp�8	�3�:L���"�pvt�O��j-��*�������ʹ��2| i~0��*̀�hQ��
z��bݵ��y���3v��p;�Q�����֠�f��c���{ p1�8}��K}���JP��g�tT0#��+d�� �Y��D�F&�b�2?�B��cm�	�Sy��??J)��RC5�vu�k��r��Y�'v�*b2^�`(��j�`�	�&�_<NP7��p�5��&3ٺ�����0p�#����'$�W�@Qc���Ƹ��8��['���#��!��p��f��E�w�^�$�C���e�6�u7{Z)�|�P��
gǢ3�\��?Ӝ��s�BO�ݥ�����>�
ɗC7`O������͞OC!��k��XEu;t�%(�ށ�UU�{xE>L���<���t6�}�F��"D6��_���EEJ�{c,;��n�bю;��2\V�ݱ@�T�����ɣ�X#yS�ISZX���)'�ج{���(���ݦ�����-��$��|>�ф7+�mk��BGi��C�5힄r49�*�YHJ�ğ��"��#;��;��U�ǚ���2n	$M�Q�8vfK7'���B�a��zh6�ʍ3J�dXr��xVf0a���k	ˬ�hSm|*�+L�����%��*g���7��6��X��ꠓh�ҋO��?zIX�0��YD��AS��=�Dw�s����!D�>��/�PV��u}C���&�>@ ;�eݵ�S���%?F��85�#�ɶ)��:� �ՉSr�*�tq���Ǌҙϳ����4�����ɜld9,��f��c���$"
JL�;
}�0�*���8Y|Lک�HuŜ���)�|]��� Z��G��rxy��t��2W�́��657ㆥV�W]���Ԧ��u/�џ�&�!�P�5������	�@��*J�`�(��B�����X+�id����H��]��qA`zЌ@J��́�� ���9�ʽ�ݗ2��j�Q.�5k���&���
R���bX���5s�kL̞֧��ŀ7Ö��Mm<_���7K!��ܟ�U�.&E�\�삈���\?'/v�Wą�ޡ<hC��}�/jp��q�6�"���c�ǑQUe�?�ڨ��Z���rv%N١t���;A@`�$�������5I0�BNU1�4��-�W�!����GH���&D����"'�"Sj:��#�c�����XXn��@�x!����L*�4��SBB��>!s�<%`v����|x���2���J��Kw����Kȩ;�!!�M+K��n���P�E�L�K��x#��G�	*��&��Ѥ�[5�R�(�OIѯ:�����$�5y11?��j�T����FL`X ��b{_�|�+�j�nP�8�t֕n7�����O���W���K������	S���`S:�\�`�t�v2���U��/����xn
�Mvլ���vA�[,R<Z|��-,�@�Ru�w�a|��}�p�2���ň���z��Q�H�}o�t�;�tE#���i���=�e�����6��'mF�?�"�%���2lt*��z�-��_(���Q#��?�e�ey���5H����:%2:Y'�������*��*'���s ���>WDI<Fj��u�+��)E����)��T�O�G��yc�e�.{��	gZ^���͓P�V�#ͫ��n��eo��bڍ�����A8S��w��O�G�a�B,�l&��d�� ��Z9��E~�[x��`r��H��g���؜"~��j8˶�]�,��A��3n�B͗^PF������X&���B6���TX�
G�t��W��6�PO�+f��3-�� �V�?����t�&�ᖒP-H��,wǷCr�!D�LM�M�E@��G���i6Ѯ7Xؤ'w��S�[�nU0��L+�&hV���r4e��/L���*#n=����,��2��3<Tk��+���(��	��\k��e�W�n7;gz9�Z'|��v]�-ilU������;29�����	}/�e>���&Xu�y���	Ǜu��Kh�w|i�K7�֝��\�G�V)�\��D�7?�}
b"�R�9BC@x5Z�˾�.ǋXϏ[q�h���x��0���-��/������D�~�IT
�̾�IJ�*X���`A;�����鮚Q��{FW�G:�p�����<�!�8g����=��c���x 3�E���J�������e�`�%Ҽ�
}^A�qK)�_��Ɛ�HA�.�Zq$X��m�+���+t5/�T �	�eߎ҄+�,�r&�.k�pP\5ʖ&�-�m�N�]o(y�~S.��DB	;�x>q�~�Q����5�e�LT�LQ*�:��JZ *D�P�p�{��-7/{����OuQs;�j*O%Z�G	^�g��N�{h�&��.>�.~GE�1��|��U$�;*����o��<�ϝ0M��[N*b�l�@6 1�_V.Sڟ`I��Bs�f�G�!wt�m��u�$;��p�Q�q�$'`�֋�'I�/�z��&�l��e	�+9��9�V���r�.F��q|zA����R�*9�hK�U,�F��y��BR�#��Y��??�Y6ׅZ��!	D��_s�3|�m&,_��0��w���4����mz6K�'5*��R���y�	�ѯmV)�'��C�e0Pr�̒�c���׏���K���E�^z�S� +;(ܢ��b�N�j����FH�=oWJE�zQl�~c��<&�K�������ͰS����hX
r�4u6c�4��Īv�Eե��iF(���bj`2���N@u"^L�ޒJb3Q���C4��(�y|C( �F���.���V�~�Y��)R����%k��{v斦���N;��q�eԻVz�r �+w�`6��J�L�a��]J�D��r_1�Oh����#ڷ�57 �6c��{HHa��`�0yߞ����P�h�8/,#G=�L"W�2�������m��"S��_�+9t ?_d�>J9��#f�p�Z�/���@���P���k\0�.��*��ghS)B:� ����=���P0�.^�]f��LW*ue��d�b�r8��?�Ķ�	�|��ݵ�`�t��\H�~,���g�� ],����Ԧ$d(7�l��
K �S�T�& ?�y�V�Y>����"Z����A�a��</�4��1�)�����Wv�0����>x؆�5�nmuǮϮ�O�t߉��L�]�~k�NQ���'��C�W��F��] 㶾v�Mp���j��XnXCW��������R�}�X<��S�r�[�$�h��
9sϼ�&��."�<��Zv�5?��kjX���H�y��7��@i���6���b����� ׊�~!��c�Z���.�����RN݊�Bjd�z�%3��`���,�q���7�M��ͭ){���肢X����:��
�#Yl��f�����"+��X��[��������j=����S1QX�eϘf�("`t�<��8�1�{�X3ob�U|J�{���xg��*�=�a� s��\c�u�ؽ���g��LY�مL�JS��%{����MD�C��Eu�%\}�r� L�z 9/XQԴ�<o�οΞ�h�,#4�Yh����G.s��h�M`rD@X{ g�ju갏�T%h<8�)��ù����E_C�p���hN�ͭ�)u��0�����N�����#���ͳlP�B�^D�p�c���#55��9ܢ��m�qM�fA!���&�/���
P5^�.����$52�!v?�w�t�B,�j#rj����E�c���_�e�p��^����!u[tt�����w��D�PD|Ё��i�Y�`�4����,�qWZ���ˋ�-���7űi��ӑ%�Vk��ϨQ.Z�A�V�E�Dh�~��;2��%�5{�\���W�6�:>y�"�ppsMj����s�����U�Q����@&�Y��A�����(E��\����P!��3JF�6���u��v�i����}TLqŦ��c���j�M��}L���ޡ W�߂�b�����'�{E�tx��T̞ϯ>:���	���y\ey|'Ɵ<	fX���p�'T�� v���*�}���Nft�+�J~��p������AD�>ߩ�f;"M+�C�0��>lgrf�R���Rr_P�VM`d]�wcӰ[���X��P�f�6�4�Fp��ಉ�g�<�nEStJT�.翔��1�(SWi-�sA������\��'�zZ�ʋ*��2U��닱�� ��VW��Ea�e?q7cc��劬����H���ٷS�҃�5�Wh��W[�'�c&��զ5R�;��#S��i����t֥�Q��|�hY����,>|`	Sh�8�q�8c�D�;� �\��9 Z�ڛ�S��D��3\:�a��GD�ߑ�k�\���Q�6|�S����C^�&�ÐH��nn+�BH���\[����u�����8�uP����oP���#�B����O?�f`���S@�r2OC�t���S�?�����M����Y��JRĽ�¢w����
� �M�祈xr1�P�gT��B�&"g'��U�s9�@� bfVvt'q�v�5?29��r�?`�B,�4{
��g:d�'���5|yoY��܎C��ϳ���ƭ���/s��P[27[ H�:!�z���FXD��ԐR _x�m�E �!��	ڳA�q�������-x�Q��w�+�76�`�l��Ƚ5���:m���q�?	�l0 ��XP'�ܤ�i
2a��[�ڝ�F&v,��Ķ��B�y�5�4�}f}1��޵=���Aظ� ���2��q�����qQP��OT\fAh)���T�֕�BG��Z`�5s
���ޮ@��^�j��J�n/���������^m�M7�P��\H��w(���{OIS��Z�+Q	��!��O���?V؂��>oA����/Db.v�?�Lj���h�E���, K���h��b�u�q@I{�a�nO�9yA�y��].\q�~�M]w�4Y�߈M�Sq� ��q��+T����(�Г��*������U��F�!!��ꥦ��h�����#�,nS���*2��]/�5Vv�I�lP'f@*/�5^Y`;���_��C�a:���`��Q�R4�o���V��?�B�n-(s���3���1�u%�m-^�U�Q
�~����9�Eѹ6��=��ї_�҅�3"��tH�Z0?���Kn�Y�\���ml�̼�vz$��-�7����{��"��Nr�T7�޳y4���bUq������"�Ak�U�F��e��؇��Z�ԧ���x��Y��)t�|^B�t�& u���6����E���,�qUR	���N�Mh��OK����x$b	�Xb=��y �ە�ɰk)
��&~�0�82`L��b�e��G�u�e��tR�J��}�4ytR�Ts�o��d�lxZ�[��}g�-�*S8D�{8���%i�.68�yWP�̵<t[����)��F9V�� ��Oc>5w�-���g��m��
YH�e>e��#n���O/�ǌ��W}}Ϫ�"��@��i�
p�Mh����1[��&B>�|�F����m&�3�j��'���E���ā���H}�
Q2?���/̦�)���?�^kh6�g��4��#ɽ��_eDzv,Ի�!����ރc�,�g�~r-��4F))�n�J��	�Z�×�˓g{���o�B53�U-Nh�{�P��S�m�S7a�=3e�ѾR�)�wI{�(~
�O���l8@O���9y_�)�+k?��{Es��f��Q�Nޞ�5���n΁Jw��Zz�uU�an�Z��mАaA=×S+�?�k������rn����.n,����r'�z���i��9�a����#��Xu:��fo]'0�ˆ
�dޡC�I�4߄}��s;���P�1ђ�ܵ�cX>T����5o���T��0�հ��3��$)�u4M`�̝��u6zp�l�$�!��g�)�.�h�}�@��`fC�g�Gp�Y֯A��%l�u��m畆���Y9c�Dfou�
���Q}qs��Z
�ch8��hl�E�U� �{�����Ƌ�v�c��	�41��kK-|��?:'7�;c|�jHt�ƪ>�P��F�{fӐ��h�mu3��WE����
�r.�I�l(���¸̘�kK�ڂ��c��4����o�X���܊ēj��&9���7?D3�^������H$l�y�x�O��k���Ќ/<�����lb@��K>����؈S�*�J���a��RJSJ�=^w�X	 ^�s��W��b��;��-P��4p�m��$����U�4֝�E�-rLA���ME�l����8��ǥ���x2�y�o���8��BI�Y�L���i��_�2M��##��:��J��A�T>Z��H�^��F�vQ���] �Чݐͪ�����j�F�m�@�L�����x���Ȑ��(���@��T����l`$ۖ���󂿠�l���!ʚ8��M!�󖉄-�=%Șq��O��b�b�"���6���gƳ8ʡ�����QÜ����{L���@�(���&�;�ۡ$36{�ݸ=ۿ\�����؎�� ���`��^�p3�h�q0&d�e�h!���w#�t��K�=��T�@�S�
\.Ğt��k�"�f%�K0�r�9��wL9��Nl�t"��z�ә�*�جe�"�:0+Q��D�6g^�� ��[#�����6��~�����%��U�Em�T�*�q҂�/��,� �7^�`�>�}����-kl����$v ����m���P�_FS*f�Y��3�dE�	aJ$۵N��&�������4�ۃ��, ������<j�������� ��j���	J�Oa��⸔�W
$�}Z"7JQ>Ϟ0e_K����CY���1�Sk+��g��޾1��O6���Z��Z	��W���%�e�A@	��4�ZTy&��oLi�>��̔M3 + ��d�֚p[j���L`N�6Wz~u6����P��M�3��#����ع�g>����y�=c��O{~9-��^�9������ng���5B��2<�03u;�\xT���2��	�|����Xl���	v��VG$y��S�N�xI�4I��zc�%'O�23�PԮ��)Y�_�xUU�je͹4��$ԙ�V�W�W+��%����!9�X��3��-�0�N���ƫ�	it�3	Y�dͯ�'�� �������j��E�̷�=8l/y��X���7�C*;kLxK�� �jҕA=��frJ���Xn�v�M]�������BP�t���]�uW�k�(c�}ک���Nb��*���5�3D�Ո/����z?�'���
.^.��ٌp�����˖��|���ڥ�a����qHL6'�%�0-Yq|��)��!���jv�g��0�̖��󜮓1	9q��N*n���b�pz�h�t���k�}/�6J��Zf�*Q�oݏ��t�r�
t/r�F�J�;w]��8y����*M�ޅMz�,�J��;�?�+��~�	</QC�W�Y{�g��� L�Y*!F�U�F���e���(�Mz�U�z󬠀��(6���D6ew�ɠ�n�q��
ێ�t}dIf����"{p>n��5��8��chG����$zcu^Ǜ��_���3�J=o�e�&��-����1���X��_��p����(?�n�Bo�)V�G��CA�n���n�"�O�=R��(m�tm޼͟�6��S��)�����<n#�:�.-𾓘r_�M�� �١yHky�@���2�3k�7�eTX��*��� 1�,�V�{��5�[�V��T�XHN��V%��wf�/"����K2b�3(.�@���e���ՙ�"x�`�3��O�DǕR�����e[�����&
&��ԥ��A�s$Y:��z%>���8���f�4�<���YW5�������DY���,�Ӗ"�O2�9�b	�O`�lJ�]}�.����2��_��8?��b	Q�Օ�����A�^��N%��9X��]+n<ÂJ�Mڭ�ab�L0�}��Z�@�ˌ��2�>^�_6k�,�#fe�\��17��N*|��~T�z��?�k�ܽ�w�3m�O)W.
������9�	^
?@���)���۬`���Ŭ�FaVo�=�/͈ШG����e2L�h�X�L�� !BX��3K�ՊO�6��u�R��|��&٣S�/��{������m_e�cʱEG8���Z����.T0c���Uzd҆�
�̀(˨�E��CSV>�h<i"X����~x3�$m��Ki��$V�us��y��j]v��,$$�pS3�X��'غY�:\38|O�-�mv.E�v�'�a��qХ| ��V���6i��m�i�s�[�hM��`�@���垛�)"X�˗`+�b"��_+$ļ�k�n	Q��� ��f �\�s'	w�b|�u����B�ce��]@�I�m���\�B}��16��C��,�`������(hN�"������!�[��j|+%�=���-ST2krXQ#�%�����69ɛJ޿ަ�q:)�:�
��i�4��bHs���eہ*�O�bŐ�]6�8*$wWmri���4�XP��!f��J԰$��^O����>����*�f�C�u�c�4����j�o�4΅.DC�ymI�ϭ�:��Z~
S�?X�m���$���Pb�~S`T��UѤ��S1�*�LI��{�L�s=�i}����ҍ��R3!=�5�&:��c��!�}��"R'�s]���2MG]eX�@d�C��.��7���k�ӯ�,�R����68�������,�wrs��"2N��튧��� ��ڊ��x��v`#m�O�GtqK�[�w `j	X}� Pk3,Lf�\9بxy9"�Ԅ:D��Ԥ^�f�.�9��v���Ӊ�����S"�c=ݠ����<��-�n]:�҇.�� ���g�;�?���&T��JV��#�P<ާZ�7u/6��(Bl�,��r�O�
�'�b�h��f{M<)E�<#)G���썠S*�g�Y�H;�6\��� 橸��}<������)��ŗ9	�_�#��]�?���32@�Ka�C�P���JuZ�ރ�GM�@�T�_n��x�u����
&��?Z�u{�-�}h�e$�9tƪ��V���k-�1%Qe�*m��+
H��􀪝�OY��[\���-�&Z���o��EE3�L�w����EK�ZG�ʘ��}�򥩅�_<|,�+��ħ��S�����lƛk��HJ䎷4�b 4Hr[J/�.��epũ��@x	/5���; ]J]c�7�,c��FE��e7�\u��5�+h����q��b;���T�������6�(�.#S��1>�^��8�a��dER*���R@h	zZu�A-�]�����!Y��<bG����;H��׮h�s� )��K,����'6�dJK�� :���|�@���XH��L�4K�v]��;!˥O��f�:�`̳$��	͜m�0r���l$L�U<v�>��[[��u�Q9�� �#!Q�t�P"�v4�+J�@ƾ3���Q�aw�._�d!�WmAbG#P X��x�)��O5��t�6디�;w*�����Y��?:��;�g`i�����*��K�5�.WL��&d�?$ 	�˳�*6T��0�9 H��z�W�v�m��!h��~��*��n"Dc�����.�)�.�U�:�w�2���"a�H��� g����@]L���ҕ�c��g �d�o��������
M����}����T����� �Q-��UZ�h��[�ּ,_J�t�t�-���-Tl�j�7��Y�nc��"_��rE]��D��ź����2t�p"3g� \C��ы"(BeF����k�5�
�n�.1�x��#N���t�����*��:�i�a����"l��*���.P��RNo�0��*]Qq�br����h���@KA���k�E��x5B�c�|��ߝ9"U@]�����+$﷛�?i�!0���X���v"�%��p�Qk<���ǘv*�jP�p����R��N:��;�.�W��N��Zxw�l��]��ƛ	p�फ़��]8�<݀ŁX� }>���Z�R�6`���`����f���ͧ�[�4c�����Oʶ�����ӤX�#�p��1�\��Uͬ�2���VT����������+Ҍ��B6��9���D`�/��"K�2N��ڌ�v�������0�#Q~��.��X(ȝ�tF�ݧ��k�&"��A�4�Hȩ�����n�����)�_x�G��;iT����WU1�j��7oE5��$7[?%]�'(��:��Z�}fr���8�X�p,���T+R��"�H���l�l�4{������A4�{e��ڵ�x�>�9"J��)?~9y��>5A`��"�~z�䫃�ߨ�Wk�3�nx�HR��W�'����򘆝ymm��Eà���y���[w#:q̼�%�����.Ō+b�3�ѝ�N<����âՌ�V֨ ���1\�> D��희�X�FlW~\0�D�u��Ew�5��SW��c�B��K��ۋh��X)v�2M\2�!l�S2��^���6�����]�rV�o�L4~�a�mkg�٭�$����֛��1Z"D�9���ʑ��:�4}H>S-ZA�hI��뛅�4��V����+HF�ءn�������~/X��9���d����çӾ{S�#��E�!4i�R�	�r�	p$���/�#��ꘋ^N�#C�"�"�*�k��GCf�=�{��Ą24-�y���~AGt�`�f(0�������=}B�������$�g��H��٘u��y2}2Y���݋ ��	pb_�Ą<�F�t��<��g�<UK����Ne�`� �J���	5��bG��kYO-��SǍz0�"<��U�̾j���J�y�H�2|�9��3Ok�Ĝl$����n�ހI)�%�Gd�Oʂ��l��`o&E[4��GM~m-��5`oVT�zb�;�ه�j���J���q����q��תU\m���R�0����@�F$Q�_�5�-��T��a�j��2��7����+0-���r/G5ǲ�Jn����۲�Z|�T4��R�OTalRuAv&	���d��L.�7b�`��z�}c��)h��Q|d�E����~�Ŏx��J#=�̌qxBb-���f�}����v	e�OL�pE�3>zЖ�bkF����[��-�3�\��3�j��X`RYȍ��o<�	+!~�h� �2výlƘ��o-���������a�2����,Y�cv=Jqqh7/Zwvu���gw�����=��A��qp캲�s�T�Z���|�>�dV�s�J}ۂ����XI4Gz�Pc�~C(a�-'l���N;I�?�]��b~/+�=����6r�L�\''�(0�0p���P�ꤦ�*�_ǲ _���f����#w�:SGچi_�ҝ�ϵ�N\����%{��Zi�k�L�}/�GA��Q6W����E��=��=�+�gU���Sd�� ]�"����fgt��mӣGr)L�W�;)b���S��v�o��G׭�f`
�^���w|���?�5���Tw�!w(��z7C��8ix��MC�� ���k���xrFB:Y�XW�`<^���������;G�G��IM�٭�]�A�q��iNP�(��a��;���RK��@wZ|��cL�ϙ������'��c 5���f����פ�FU�:Alm�I
�k����%])٭�J��㨨nЋ���¢j�
O�[�q��s4n�!�YD�OZ���T)��������z]�����S7�ׄz~C�-Y���NN���!�]��JWх�B�u�9��P'�\4I/�^�
h���J���#�8@q�܁��G��1�u�S�6����H�5n��p��L�W������d��\ߕ�_/=U��th'1z6�0�v̲��Ǣ#�ah�h�Z�<�����í�rC5-T���2�ܱ���$��ZU3
�i7��ܴ�H�8I�q%�z�����������=����TًZ������qdj~zo��}��(f��|�d̞%�Φ�C�3��^xN�C���3t�"�;T�r3h��.+;ع�*��9�|����,�D�Җ)�Xf���+�q��#�$t'I�hm���oc�ozxs!ߋ�w�q?�?��,�}b�E��$=�l,_wif�� 32�-f��L�.h��/���Lj'����a���눖��
�A��{��S��12��/3��!�}w���tq��@0�D+��@��/���886�(�`Ox�S����
y�g�����q���\Gu���S��2g��{S�����3�v�}%�E������9T�#���o�Z�����/��x�Y}���D<%����;��� ���lQؤ慄�4�Cj���pq`~+q�Q��%X��RF��s��"�-���C��TM���=Xd,H�h�gp���Z12�YL}�ᵺ�T|�O4�R�gZ�8�&��?����+2���ã��w�,<����è�#�Am�̲UY�L �����țl��`�'$����N��s5�gp�ݒ�jiӚ�J���tA�a�W�֥ :D��j�ٰ"��y�c���:���&��Z��Tv0eG� ��[��x��w,��^?�He�T,����ɳ���MF�OM��`�EK�?�‡14ʩՈ;|RȰ}����הW���B�-n�����[�}q[�m�zda��~�	�86m���_
_N�xǳO����"�c�;�,#�Q���6%yZ���Hl�eD>�e//�0{el���'�<��<"��yB��<yČ@�:o~�MZ2]��2�7H0H�z�<� �S�ĝW����}����,=���K$�тъ������5�eN�<	Wx�u1Ӿh�6w%�}��I'sk�2ըިR^�pZ�x�H)ɺI���ڝ�ubQM�%:5����!��]
�Y�	������0�8$�`���u"�%�yBOw��j�2�r��_�Q{�^����d��zNG�����d�=Z�����z&���3��������y��u��d���R�',��(�+���̛֧O���P- �t4����:g1��hWu�ˏ+���J�� 7�z}X�N\Q>W�-�u]�r�sֹ�&ɳ�-k�lY�B�}��[�xm}H�_�#����,��;HE����;�Ώ��Oh��Zh�w֪q��n)�6Gl7������jh�{�;l_��6@_̪C5�c��^¾n���D�]iǥ�Vdj) �.�� �W�|Ppha�X����d)�8����ۀ�S��F�y��m!b��ӓyg�R�A!�V�_�s�'eM�I6W�ހM)���������ؚk����:�NJ�xk� ��fX��D�"�:���B5b�1ߑ7=
��ЭNU�%f�h\���7r�sRpU�|!�#���pS��H?7fo?�04f��e!C��Y�G��2�Q%���#�C(`ow+������|l�5�;A�5�A�=~�Â��*1耓����C��j�uF�"\Lܼ��$V�Q�u6*�,���#�{������yW+@�+D��M+4���zy|fėvF׿J�Ȍ$�gB��u �Z��҄!BK��<ٔ�5�#�p���x5��KVNE ��@��yz�!#�պ�Sj���V�-�����\zkք����uJ��?	j@R���a���^I�p��Gi�������rd��٬˻��_2�[C5x�.LL�Gd[���kβ�	 S�ƣ�d����Ћ1�үU�&��ԴBR�+��7k�G���L��H��`*���W|��U{~ �8���-�W�\,~��\���qG=�B|;�9L*\ݔGg]��kDۋ��R��u,f+�����d]X��y/8��R!��X`�@�A^ՅP J�
ɓ�E�ě܊���J��!.4����k��`�'5@��Z� ��U��*�rrIO�sہ�HG��g@�c�����
L $)�s}ӄ�u�<�ؑ_I#�g���+�B�*�Q�I��U�2�t�0���Ñx;�q��'��{��Vi�������>0��{c�e�%�7�!~ z��������A �	��0k���J·��(ݬ����f���/�=��d
b�~B_�x1K|:���|�ߧ"�_")�*=$��������D"��hr��5V�����*�#�M2ӏ���ekͯ:���� -lkzI�$ו��0�I&�8���z���lhď�c9�;"u��I4��_�"�
��_����)B��F�)�cu��y�Fn���L�{��3�z�d�����h�	+J7Q�X��BtW�,q%��S(i�)��L�n��GҜ�Xv�l`4�-`�zbD��O�2+�p5��_��O��Z����ڹV�ж��3Æ*ۜ��۾ʥڙ�R*���!+F��{�ZWv%rF�D���I��#퇥�m�%��>�����>�Z���y"�����aW��!��U��:��!�bm�aE\�`2G��CFf������y��RLe��e���CQ���6�}�KPN292�ܮP� b�	2�� ]����E�IN���);����͔� �����+���s.�̾sH;�Qc7ZՐe��׍:��sA��Qy�A�Ap��V$d�������l��c�\{��ڦ�Q�6+I���8.�#݆)@���U��a^�_��4Cj�]���x:x�JC�1��'O��zeRP	|��et�/�>Õ�����H���S{�,v2��y]����MQ�?p[����8�~vG�,ǩ�F�&�ĄE�p;A$q�L�9�^cŽ<_�,+��g��*hs�����z4<b�?7��E��o��e,��0��{�x]@���AV_����=d8,#h����F5��
�Lݭd�����n��5��&>܍� �}���i��4�1%S�
�x�u:�Z�FB ��,&2
hk��Ɣ#����m�y�c�?ʣZ���@wI'���@��\���š4)�X�k���e��\��n�(�b��N}�ָܪ�H���t벜�p����H�)�qyYmif����#R�cN�J���M��4W����y��&3>K��kWS�8.-�=�
�������B�Dv�`��Ksœ�� r�?&��U�Op�Ӫ_�ֵ�����OX\�Q����B��3��\�h��|��]�7,S�Y�?��^�
�V��Ԏ�S��:^S�ࡁ�w��x���w]J�M.�..V���@�ĩ�߸���-����P���&��vO�g&��A췢�FM�#1HT�F��.r,�Sa7�ھ� �h��r=h*�,.�?셔�u���X�uo��E���R^�1�ˍ*W����yZA���,����cY�oE�@�9&�
�غ|�0Q�<a�8{��Wק�
^vR�5 3���լ�%�>`��Zi�6�L����<v��*X���=����}/�ҕ4��|��fS�$ZՃ� �p�
cB=�	�����>N=ۮ�c�^h[¡t����v��������7%����18G#���8��v41�6?���T���o�
���_3
Ml5R�HnY�S�GG�,欓6Κ�&QJ�/�O��s��dx�ID@|Q � >2�祁��<x�za�C[��(�K0�|E�j'�H�C[(p˕�=�[~���guG���2/E�A�C?�?�b8�����=���h#��,��)}˂.�Y���ۚ�� �ߩ§��9H۶\A��r�yF����by�{]#�X�͏M�"����KG�%VM�@�	�j���z��\jz�#���C�T�}��y�Cs��R{W"�	�{�r�\�M ���E���<Fv��+ԸߖBq�P�Q+ܲh�/4�n�O3c�ۤ�G�z�����)�J����5E��a�V��hҘ��hAM�c�wu��2�Dqt�#
�Lֈ�*B��/랏��߲�S������,�L� ������/{0���h�2]	o"�ǔ�3/�^o1T�*v�]�Qcӥ��������c&�r�K���xh^�%\�V��$������t�R_%s�q;TS�_�Z��ݞ=�Њ'D����.��S�(!�3#z�dj�{�6�犡=8��-�C*C���Hg��K
ё����q���ljT���Ԇ���.�I��<,x��r���62���1�˱���Ҋ�%1p//_Я?M��H<u��U��J�&q�0S[KIQ�w���ؐ�4�7D��
�k<�"�"@?:OZw����i�=7�]-����
GZ��@`p��������\�d�Q�న�V�����`ڗX���J��8��A�Eak��Ź.5G=7���Mm�^�T[�`읤̉މs8������P���I��b&[RՏ�W��F9��ODɞߒ�����s���B�{J��׼�"RnJQriT���d"Nj�w�4��d�)�x�x����tw{�U7�˩$; 4�["6Ƅg�7�n(E"��Y[�g�í�i��xR�L�W'U��]��b�����FQv�x�Ok��\ar�1�*�;�"�6�i��ܾ�l��srC�/D�|1K
�5P*�V�?�Mk��PU�\�@C�12V��D����WB�e�z����z ����%J���%R�,���eE��E�Z��	,>�0.n!�нV�H�T��s#I/0~Ӕ�@���܂́MT�I��`,����r�\��u���D��u�����s�
��8�/���-^��F��\V����-�|M;��Mp�[��T8%�	vy�u��%*��M@鍵$��&�0w��S��
�޺uBr�Q����&֋+D���Y���ر�Q�z5�6��k��4�bG��X��Hmу���~�z��d_�n+�(B3|��V�������8���I��=-:*q����6X���MII������~VT�z,N?M���/�N�0 ����{��5=��`@Ԏ�����yq��gز>�µ�Zr��K��F���_Y�L��/���o��ԭ���B��r􈒇�x6LJǇ�Q�r3�h�0�2f�As�uݨS|C��7�_�h��6��@�[8KP#ur�v�C�e����Zz)#�-d�$L�J����5�5(����7.|l����Xi��yӆ���v_��i1��H���>��Đ���R�E8��!��6��2���M9-h��00����Fi�h��׀���3��ʥЍ�p��F(�x�9|�b*�"l/�Y��?���r��j���7�r��H4��<<��
"��pOPW��c��zV!%˿�\ !�|Qh�[��ɲ�:3�C����q���|a��U����wD�T��£�,"Bs��p���G���zg�Z�9���SՎ�i��P����Ձm3��ZU�R�,�Dd��$�8!�}R�z�G���!�9��8�-[!��+(��}�B�;���	Dة�]뻄�z�*������j��f�I.�ьL0�{~]�!҉�z��J�:�S>��6:M�f���k�5�.E��1�bGI�F"����7q�!�WN��Yfu�juΞ�l�@�Ļ`���^ϣEbwS
���$Ҫ�ga���_U�iYR�P��>��S���
ZG�,��ȏ���܊W�3_U�����o	�`u����������2Kr0�H)�P/�_�*�*h��Bs�(�,.q	�G�9�i�^u�XcO���r���&�MkEQ<��H���x�C�ERpJ'��@7�����CIZ>Yݤ��,F�lE���8�����e�p�:z���$v�p��(Sq+#*_�#��z�/l�޼�ƣ���ַ��72��\�՗�q��3����}�D�����[tl�/�0�Y�L-�UM�����/$���k�?����'.9��Z�s�u����҆WxVW`g.�����y D6w(��ˊ��O�L�	.���I��*?������0ͺFݩC��p�3�)�b����i����A��c��r��r��;�G ���ޥ��N��0tW�J�4��F���̆�Z?��0������a��0{Q���Y��
Y�c�*�r@z��o��9M�n�J6�4�]E����B�x����&�w*�#�����Kr.Ъs!��PD����5#&�S=ִ���9�Ob��A,��L��c/���g���l�M�|� o�o/ja��TlYm<#���wH!6��h�+^�S�tY hC�G�8�K�{��6�]�&,���J�i|�z�d�f?*u��p��+��l-�F�M3{UׅY�Ae;�|�$��%�t�@�+��1G�z�\�u�����< VA><c�"]D�1+t��Z"O�����Q�:R!-]�״���r9Һ���Bn!�&�������W:M��q���t+#a(�F<�7�u+��;��|��쫺|�2Z�-�7r���r�ZٿFF�~���ٻ���~/,�0��WP��+��H����/ȡC�染,ZWi���Yb�*쿳|��2��:'˭����j�1̞���|+�#�B�EOF�2^~"�灭�>��rI���x���Xr8��<�W�#�ޡ5-_�8	��"�te�M�
pI��_y�3D�E�ӝ�]���֥VZ��E$N{�Z��ƌԱ��^��i�B�s�ߦ�ty,��Z���&s�@y9)wSϽN�4Ĥ�7H�ɻ�+�<`lR� `�zjfw2QƗd�聰�P_]>E:�G%.�-����<&ے�b~�Qx�����o4Q���XQm�9s�����q��'xy#��Ӆw�¶.f���G���q�]�k\X�j���(�o�~��b��;�D���3V|ޅghb���u��Bz���H�$��I�׀�X�u%�{��((���4S�{����0�n̖�u�j�_��}o*G��K�r=�R�Zz��|��h1��\��e3�p*��K��I\��.L9���Y��z#�pͮ�.ZI�
C_G=�6GI�\�{��!�����5�MvK�PJS͐*S�#�2h��\����W����e��k���p6��3�_��ҭ��a��q�\���'36�{�A!��&A�`~��~>Z�qC§f�l�+B�'=�R�=��f�i�n�)u�������oZ��a�-T��\
�����#,�ηw����f��#��y�7�^��#��c�#H�މ%#�6%��5���������9�݌��<R��L<]�,�X@x�~x1� �� 	��-d���U��\��T`8��%?w����1�u�n�8�q��!��C�n�n0�C&Ѹb�e�0�T�Y�[�գ !�3�,����г�: ����դug�0�� G	�,�t�N�o�!������t�b�P��rꟇ�DZVƊ`�c�e/�v���FC�,$ъ OIQLd5��͊_��>��\wk�����)p-��q?�D�Z�v@�!ӓͣ��I�ثS�hp�L7�=Y �����R��Z#�����Y������5`t�+(��<C��1A��
u埭�k��l���%/ʇ�����a(g��G���P��6"�6OW�јǚ���K�XJK����z�����^,֫lL��v�	v�-�#���Qd[�(�/��#bf��6z���؏�h��{��R�uUkNR%�o�y�q�a1g������4�g� ���ͨ�*���h��z��K���eP�I�y����l�~�6�!��o�lt<���d㥍�U�?�[5��R`��F���L�ek���pկK*�+	��#��7��$_j���d���4Y��{�U�/nR����(�������'G.��}����@V�2�C�,N��k�4�O�7mǭ��_���f~Zd��nu���M�|Y�F�kb�Eq�s���M�	�=�a�jOH﷓7���43�������b��$v}�S@�sK� Zţ��2&�sG���2A`�c�X �Q��'��R�r�)���,���C��+�20/B��,FLLj8���+qf皡7&�hZ�y)��H�� 6#���k�J�����嚉�R��t�����%K�G�6*�|�izj4a]_'�VѰ�(���)���&�Z��=N[��/������[t�
1�
�[�:���'����d�"��'?a=X�}hx�:�W�;Ԫ1���%_�讠�vikT�D�����oN5`�h�)�Y-h�.��� %���Ԇ�4��Y�LG��;���������Z �f��zl��<���|������V���n��o����D|B�.	T�!�P誜[�n�J��c��b�O"E�Vi7�THg�G�ZA+̺�s�;X���%	:>jŖ���@,v��ٞpr^Lw����F��T�Q�����m��y��]�#�Ǣ�Ҙ/i(�\�P�_��Ln���Ь�
&&�@瞯�_O����
��E�mi���;�����DS���ٲT����@�g�w0���TK�Z������Os�ׅ".���WQ~����l⅑���6��\�Ų�lCD��@b�7x.�6
�&Ϟ�	lO�8��c��+����a {%��^�x��<�0<�xG�q?�nЦy��v�^����i]�삎�`G(�F����E'���\��e��$�>=�S�l T�UǇ��	7?G��/�e�\�����Sc-{�s,�M��~>���c�e�\�����|����r��%/tD�e�O+�dج$ @S�w��wͣPd��1��N��Y�6�YUf�������L�S>k�:~��:H�
ɽz��O;+��CE�H�"t�.۬�˔R��Bᣖ��@G�����k�=�%��BQ`⡐��/�gӥVԡ7݃�S.�od���,����=d�G�GS���g����������C;_��#��`�3]�m��ʦ�~ޓvz�L��<5��)Ή��`l�� Q�̆�0����Cl�@���L��U�6���B�z��s&y]��D.�[z�� ���p�ޙ`�/xȻ�!�f*��8d�D[Lt��4o�`���P`��r�tuؚCc�+��kLi� w��\�M���E������-酇��\�oF+ *��wtpqB�N��:9������'ڰ�LbL��1N���)����v�A~��Y�ƞ�]����;d�����Ŭ���Ղ�'��M%ƛ8�{n�:�ݢl�.TK�an�Y�:�9f�m	T���Ud�8��I�H������"�Yr�4�+`��cJ�PJ�L9���艽=��Z��o���s��fS�d_�E����̰%�+���p���P�mu� �8G'�Nz�7�0�g�i�B-�U�]H�iLk�c�/���u�������W���)��$?*�+�tG�1�5�B�vY��H��PW������%ߨ���Ҟ�r��vu&�bg���������*z`�s @=o��$�sQsOp��k�9Ʀ���zl���
j&?	�H���8
�s���2Ghiy���L�}
�jB �i��݇͛ ϱ9��TgǢh+�e�� ��m���1{��{į@'j2B�-���F�j`es�%����� \�,����]�;u�`�	"%a-�>ޯZ�N������ ���f_�(�Ǯ)�+��[I�V���2h��JP�e�13�m�&��F)�(u�9��{��&�?q�<Pˠ�o9��It?�qg`*zD�͕s��DU`N�2*Q�&�z6��������pwy���*�0q�m���JP���p��$ϲİ�vb���\@���Z�����9bՃ�6���\(*�9$p�"��{u`��ߤa��β]�e�LC�9���*� ����* L$�4�e�R�q{E���C��<�)�B�����vV����	��ٜ׋x;CKэ�5��f%��"î\��EK2��m�k�`��E	Ϋ;�uiy/ҡErr[(����|ms�۠�K�8�#n�:��8��8�1z��
�g��P��<WB������N&C�Y쉒���1������
�痽��6�N93@a5�t��.�T���)���-74x:W�ȝG'��}i��"{N,�I�e;T'���	�(f	�	�g=>J>�b&��b��h��'�r9"��������l���R�i��|���.�;���#!$� �NUwSj�X=j��
(P�F�;���E�E���2\Ic��V�E�I+
6�����|I�JG~�w��T��5�al����]��^G �)�_�Y����[d;�C��Td��U���P�Ŏ�5���Ea���f�J�T3�v��p��k�́���j
m�z#^��8=��"Č�Zx�Hf`$����ӎ�P�$����<�psS�ReF���4�j<Ƚ��Z�ܹ�c?R]��L��{1���Eb����\����*t��:�巒L�k�ԣ�[ �2�2�1O�����,��k�4��7����5�bd&�٢(f�d�A�z������"��w4�)��Ϳ���܉!(����nV�%��}���?��I7w�oYj�4�\]�&�]����H����js��[S�+���t�؟F�������[K}�
���)�<q���XVL�߷�EMg�d�[�AF:�������s�!�;������B.c����X,���7Rz!�{�5�P���W��}�"�y�0A�HjX��+-nG��J�Fxh{'�u=_7ΐ�Xui�52n�ݙ�*#�L��t�é�#W�'Ը��1����������ވh��I[-������h�g�3���G�8|3�87�)�oǌo=�+�,W�
����2��f��
��l��ۣK�����˪��.Ѐ�|k�������fM��~�vO�ŏ����PbY/Y�05��o�n�k��|�u���E
�n�_5L�jru�����I��z�U���M��k;�r���L0a9�(�-6�R�*��V~4#�pa�T��N�E�\��� �����݈��O�D��ءM|5V A�N������mC����� ��b/���������}T�6�ѿ����s��^�&�nA�ԝ��?W�?��O�c�Q���q˷�u�R�'7b_��hu�2>�e0�H՝��3�D��5�!8�H�L̓��:��p�A)L ��7� �+����ƞ0��V�v��,�8�/��2�_�4Y�ڤd�yO_:gv����*���%�^���W��hB'��p�d����n�k��p����̋ɄD�>��e_Og{�\Z0�Ν��1��.*������}r`*�z��\#�Z��i�S�i�6�7j{Nj�D��g"�j�Yοtk������+ջ�)��៮���+gCx�=������`>��c��)��۪��-~^��H���bF��%�$�
�,?���+9�)4���.#ͩ���X`:�Z�`�����l��K��x�����`V��J��x����{1�^�<���s��Dt7�n�*��Hc8י^�(,2O���^997CXL��2�ΰ��ƝZ ��[rXq�Q4	�!^�Eu���fw1r�t�1SB~�8ߑ_[Y+2�ߟ���Q��Z9N��;�{��(ł�g������%E����i��s� ��"n��}"Zǀ[S��l^��ƈ�l�4ܤ0{�$-�7K����v���-��gx2}mlX�:9)~:W (Y{˝ĳ8��EpZp*[�T�`�!�G�x^�[�x��CX;���vJ��xѳ�ʓ��{�SFͼ�4W�s���\��R��;,�GaƮ�{ ����`Q��e#�BL�f��qI
��)r��O���k�#�:um»�^c��T�7\Ȏ�V,��L�[T�UG>��V��g��pj�҈i�5�WΒ����͛vF�-V��A��M-��~`\��&�D�ih���Si��e̴;] �ftF��t�,�I0ʣ���:J�;͈K�J�������A5�����(qr�Dȧ�O��������r������ӂ��'W̢�$X��^q�f!�(��ƣ�n �e�4�D�*�0� �S��c�l3�	H=X�>	f 6�ƹT��M���*=�Xyg;,���p�Rf�i��������������1N���$��9��v܏��k���I�1c�[�ђ��3v��ih=��@�
�j��^�����#�K�)�1�+�HhU�U�f�%�*���l�Z�'�^x���?aw(��vL	��:*����k'�P������@�!uFEzb�cT�1��p�A���M�Y�WE<��tC�0Ǆ`_��iL�j_TiЩ6])�)��D��C���X��j�����HKJA�g1����yH��j3#�c,_"��7��)0�_yI��H��aJ�\5;bq�p�����-t&ί[hXxs3M	��I��Il6Yf�����Rs�w��2x�U7X��OJ�t�z��;�6g���Wb�/[(��_�a���]�Д�9����&��������{D\�(O����hI���s|�w?:#�t�	a��A�)�����F9 ��e�K�3@�bʢ�JT�m3��F��R�7���,$���9��nf�N��W�N��l@$�AV�����B�q��VI87��6�������#ؠ���`��L�[�BDZ�r�b�,��g;8eϢ��F����[�J[��'L�ef*��
G0Gٶ�cmYzr�d��A��zr}�.����J2͠t��Z���Vyq�M�e;6�����e�MZ��;���_�ʘag��c�����w��{������iA����������$���OhnR��ZnYQ��A;+N�;ǂ�nx1x�a�V8��ן��R��<��������	�M_�:�p����P2����d1����&��5��[hI��X���6w?�"�����s���	��>ģ�w[��xAۚ���Ƭى�2F�@��"�:}�&<aBp�P<0����*����g..)���6�1�FE��߰��/��Y����x��<�~�� ���4a-�:�4gO�|"ymkk*	O�����������#�.IsZ�B��.>ī�@��z%�x���%�+X��I��i�-�7�!�6
�ԮW�Ө'ʡ����n�����\Er[��d!ǽ�hI%����� �]��'1jj�O�J���G~G���]88л����(U��-_��4`�{�|���p�X�P�t5���F��գUԐ~
^��\nA2+���� s�Njtj�+��e8}0sVQ�����-«�II�2:�=��k��F���D�e���]���oA�j��|)]��L����J�f�E?ڛw��f�!�Wދ�ɡU\ �;�iw���B.bYU`m3�6���N"�`�l50�j�f�~�l�
̍�@�d�'Ω��*�G��M��	��5GG�Z֦���pn�\b�� .��>ң��ѣ�zZ�������&��HLq?�f8�aǥ	�+�A��T�[��<�G{m�s�J��v+����VE=KJ��>��&���L"k�����Q��A`�G��	@D]�1�P/�z	�%�z��Xk����Z���w�'�}h�E��\�HZ�E\fe�aD�2%�f�5 ��A�Ϥ�>����0ѴY�k9���V(�=�SFЦ���1��H�ܧnKݔ��N�oވg�����"*ؖ�",W�n}�n�<�-�����tL1�zE0����O)l5��E��>�i��+qI�{
�_��**S���~l����q56�$	���X��Qz��.Ʃ�N�|U�������+�	�׳U�t΋-��VH�|�p��S� ���RMֱ@k�pK���	�iO�:��"m$��;��)���\?3b�l`��Y�Ro��C��@�9����)�;���A{0��*�|���a�-�ݸW��u�fuF}ƥ|X��R�1�F&f���s�����S��כ�F�H�Wg[�����Y����j8�nю$�F� i�RHf��J��6�j`1��g�i��N��"L�Dq�Y ؚ���A�<�i�S�E�r��hb�.sP(3XU!�L�2���P�@��wt��b= ���w؞����K� һ�D*�<�/>�B�am�Qw��j=�&���D+�!P��'f;���
S�[�G������֙�Z�w!#�Gԟ�K�����7���\,R��-�[�u�~&�]�&8�ضF�	pZNX|�m����p3��t�I�w�xr�����h抇��mh�$�#Լ(��o���7���	�TL�jv$l��Jl�q��r�y�%�H=R�"��X��,�!h�So`B���Q�an�c�<V���N���xwt�ĳOm�sIF��̷_Ʋ�l=�A��~�ؙ��|3����
v�/DVM�<����!���+������L޾r����;�>�1����O��u9=�.��uzˍ���G�o����'��iA���o�Pnb�D[�cF_�Ler���e�x�����N���\vj;3sH7�U�w��*Qb*��q�Q�v~�o����3T�XhU��j4��[4��
���l�!A�zťq�^�_j𮫔g��dc��Hg�ĥ`�|}��e�
l@��Wp�.�;��&>�y@�����F5��n��P+P��#>�ݸ%s�M�^��b%K��>��h[2�ߍ��C��Z�f�ڟ�f�~G'�i(E��h��JſU���/�Q��ߏ�z�'>�j�zI]�D��1>�/��(���K�B9��U@d���^���Q#����MD����K!�c�-�����e5$ܡbdz0/�7�����Z �I=��/�UeУ��γUmy�I����וG�P���5�HHm�ߛ�t����X�����Jw`��in@�dD-�G��$a���>��Q�yiiR�ͷ���b���/���1��irW�#�ƿ�q��P|���g<��3S-ݐ�	��<��zP�q{����������{	!�]������ՐC�ֈ���1xG>��cE�nh"R�2c����^N�l�B��4̣�wS[]�����jr�g%ĩ8Y��V�6�ٍzMU�֞�ێ���rwo�2�E�j'���(h���v�k1bw�d��	q�j��[ 
�"w�_��5���A��	6|�`���<Kg�([L�ov*aC��t�V�MN�w���X�(̂<b{�a�éH���F*C� ��쒙cG��#��c4��k=�=/�4$�d�P>��-e���ԋ��������j2�!`As�dT��cP1C����,L8᠍L��[XA�z�#�6����0�,b�^�7�P��B]'[�ү'>���w���)�;G���VXI��]�R����k{�]NH���Ζ���L|��#5��j"�����P���t��'lb6��Nڐ���������2�������o���PHN��e��ۃ�F���U�_�❞#��Cj0Yu���S�"�����
h�)�TD�UR՜���R��vKH�6	C�b����x�$q0�����SX��M��̆�J��+(��<ˠ��W��О98i��:^��M��I��k�M�(��5^�/���w[�R~F6���-�S�A�>�ԉZkQ��g�Ӧ��%�J$����S���U��)���+�^����v���[�����%�G���F���X:뱗z����g�p��=�$zӺ�����/��B�bh3��L!Z�Uf���	��t�t�z;���e������^/�M�h:öb�K�?��o�̓��6V�i�� ���>(! �|6J`C�����NcF�lx����T�C�u�3�a�{�Ǚ &����d����WLE�Mwɹ��/�Qw|�s��7|�l/�^�=܍aj[(81�aB�+&k�,�< �\W��NP���A�=|gx\Ow?�QݰDj+PN"VX��^,�ph�ϙ%[�r�~���B�k���7i��,�fh\�C�gO�qi<��L{ WO�$��g����S.1�sv>�"u��ꉆ�ΞI�<�����>2G�0w��x�k	��;�"q6��Ӹ��i�ݹ%��4u�d����ڋ���䌎�䗬����E�۩���%(1?S�����@!���'G�«CL�C�1b^�G���o+�����R8GVMA�.,�h��"�Se�0�ί|f��1����@	�ڈ������"�'���H�����$�[S�(�����@�����a��ՀI�1�VZz�ۤ8�Ź��7�:��d�shv�B��_K ��T�I6�ě1�ˎ>to��ww�m��F�)$ڌ����<NϽ�.�b%�ȵe�`�n�� ��4�� ٽw,I�T�+��&�N[�>C^8�C�
{��x�f k$��j�I��c*�;��o��Nf&��Ԉ�ܣ)�@�m)�13��"Nl �$��ʾș�:;��7��G��\�bE+_��^x��d��2c��8;�̫��]�n9dB��i�_�E�>�����[�:y������Ok����C��^��lW6T���R�Y�%@?v��Q��a�ܶ�k>��Cj�>7���Z���:�z�{���-���zv/E�K�0��p>����n�p>�����(yMK+I]7�@��W���Րb����HЋ�r�E��fI.;Ff՗z��"�c��L9��X-˅�C蕔�C6�o�&�� ��l̰l��ho�K�ПA��siK`�L�ÒT.�+0N��5�SڣL����$���-��UV������v{��=nc��N&�	�� ���U��G�T�KĀJgc�P�#~��W�n�g#�����t�5TY��W��P�����l���]i�W��1��"o����������"��j��
���n+�9�m���>i�@����0�S���fC���3�k��a#���s���&�B�gT���}�������'��%���Y�3	��p�PӮ*:	RJ���]q�r�N�&|ISC��\�����E��0��7��(-�5�V!W�M� 掣�c���~���<(�C����+3�' �:�+G ��P ��Q�^V�e-FW����3O���ے��������1ҹ,2�/p���)���p�a���&�f\��pUb�7��N�����(����%C:Ƌx��)?�D-�*��7���pT;!��}���V~L~Щ��/��i~
V����hr�b��ѩ/�T���QMԿ��S�I'�w�,� ��\�8�)�ꇳ�rφ��`%U�]����/�35r�Q��������xS�n���M��w�:fjIi�T�-G��Q��{���|�K�!�xI��Z��x[�@����b
��GXI��ħ�1���z	Y�е��^z����?���7���l���y:�� R�;��ׄ��4��n�1�?|�^S�0�̥�-���xK�j}�Cs/7��MUρ�������� ����͵�mk�,��`!zh:����mX��#�q:HA��K+�&�]^�ΕÉ;߫����&c:f��� ����,��h
�нT���qw�CL��/F��v�}��,eb'|���ܜl���Z��Ȗ=^��� �����Ѣ�\\+�1��$o���.�r߮�(OO�>��v
�D�� �� �l�m�WD?�t�%Ĺ�i�����<��]��r���#�}Ro���q׼�ǰ'm�鏳!6� �]#x�$c���B��A����(9d�6� '[��pbn\tuw7?��y�|�X�'��[������1�[ny�i�,J����K�:3]�]��^x�w�0Jk���a}�a��Rn�n[�����bE���L�q�K��ֱߋ�F;79���֛�u�B�g�#M ��B��-�T�/4l��w��D}�0Tf��tÀ	�����ً��-�JxP��ܷ쯂U���&y`tl�хV)zC'pck�_8��Y�P��팋���*�}�^-�浏����܀&Cd�x���uS���)NL���)����J=EUx�8��Tiƺ�ڹ��}�ZG|��He�x��^t(�:{<�XUޖ�-0��F���*}�,�����ގ���M��=�A����L	�X�=��`y�g���?��P�Y
��\hNp�9~,W�ѿ����������D�2�0���Q+X|n.��9�8���aE��s�(�/wr2��|�զC��o�"I{�G�A��.o��8�˭���I^*|����=�{>�Di������0������1����H��%�7g]晡XC�:����c�Y����&\� ���BpF���MګK��F�ik�����7{3�g�4RՐ�A�2�N�3:^�E/EX`�]3*%R�x8������@�J|zS����� }���b#ޤ�C����I��5*�&�(�2՛	����+l{�GA�()Ǆ?���4�/lJU~l!��J��͙��q�)8e���s0��� nr�9�Y��k!"���/-��V�͕'7d�_-��+�0�C�:��2�Jg@bs�R�f����T�|�������i�W�Y�P�r����X�ב�0@Z��Yy�#ZVG�N)vI����G�fo�ucy\��բ�;��fr:j�jQO�#厚;���Ƕ V��9�=k�5>����5?uuP����C�>z�H~�;����Ɗ��90$������F!�EYT�@�(Y��{wѪ���R2�!�V(9!ޱ�`���m���Tf�'�	G���P`ce{	���B5������5�d�SG�g\��S	�d0��D��2I��8�!��ƛ�J�""�V��� ��a�#���T��X<.H#�l��x���t������n.�>h���b�fp(���p���#kl�ԌՋ�|ΒY��?�c�Ȧd�z����l�S@��BNw�Xb>��]s��"W�S�Պ�c����~L^O��YNڠ�?�����"�6�y.C�[rwk���.���}ɴ{�x�'�e��u�4r�#���)�=���S_肠��ިKV�k�L>ߑv�,����6�|���e��Y�{V#	��.��D���ն��.ڦg���G�������$�xŐ�w�s |��V�XՖ��y��v���\���.�`|�M�;Y�7�ko��E�	 ���r�%��ʚ����@	S�	d#Y���H��߬yb,�gI�R*I�QEB�u`�R��a.:2�Xb�첵�����ړ�*����m���Y/����e+�TS��}�:��"ȝ��N�B����0�-f���ȗ#K�	 �J��K�
ɿ�kԖ�4�s���Q��&6��(� gP�/�O�Z7��fp^��τӂ=�3�pq�n��`,��+.�A烳�cq3�ӕ���-lޒD��Yp�]z�Ahf��4��̆�>w�z B.kI��Ėq���j���|L��_n����}�Q!�����F��4�Bp�=�Z}^�x��.���S/�	\�X�➸���P,L��#n)�ӈ��\
�^%�	�<����j�n�����1��)&.%�*��t��}�zJA4�N�-�j�1�s��ڬ�8�V��$釉w��|�X_�Y	ilMj����/+D�b��$�b>��juH�[����l���e��\�'���~����
1C��m��eu2V�jq�X%B�Y��9	d���sj1H^�p܇�	��-
d[C�Q�xM���/;�A)Ӌ7�'�ψ"VH'?�<�wHy��T+
�Z�?;Y��XT��h�F�NPӋ��=.��5�¶_��]�=�����쬴x_D�Sw��c���b/�����E����w2��3ϧ�\���.�wf5��?n^�R���<BKW~%͞ɛv1���ɬ�-ke�6�ܿ��ri��$1'�$t������`��^N��)�V�g���X f�����VJ��/�b�8��4�ɣ���)SŪ��٤h7�pޣ��+Ѥ2�_�&��QM.͒b1�ςS��|NO�d��mkWzuzo!i��.���7F���bB���P����]��D�Ӿ�,��6�E������i�ڰi3f��1_aN��ՇU�E8�0�W� �������!�_)(�t�O��F��?�#�7;�G�]�>�ɪs�Y�$e~:�����)5��� ��L9�ڱ#ђU�@��o������a8a�0cwl�A�݆�%��}�F�MH�3�-��U&B��1��)�˨
���|���]v��^�Q;�XAV�������i�Lȝx��!��G����ӏj,�.6���:9���#|�L�x��SA�5l�P�<��s�G¢�����Y�5��Le�;�T`?q蚙�Z���6>�pk?��!���{�����ܤ�5��$�}V'H����)�Ϥ�]*#����c��"g���|qf*Pf{�zEr2���W�w`w��-#��δ'���N-�����w��{VU��CW��L���!7Z�o]tˊ�j�=A�
�q��]krd�b�=������o�e�r�U�ʁ�=<~X됆�����syH�V��5����̸A�ͶQ�wO��z��c��G����Q�-�&p$}"F�����\U�==��R=�AE����ϊ��K��ĩ^͋0�m.�u�jsfʳm�ƒ %�ؔ��T�ԥ�H���v�:+x>y9��Ut8@����?���O"X��j|�U=6-���u�8�^�l҄�m�Y
{%��&o�5��e�N�5�Lb;f� �n����L�T����x�l�o�\��G�
��	��v�s3����o���?�y�J�x��j�|޺�B�V��Ts���D��-:�O@�"�kH@WN�7���X.��Z����$����eDY��̺��� .�05�|	���j-��r��^�I��u�ā�P���a�fV.}�aMW�=��t�N��;����kH��xyI��U����;��b^�~4y�gR/bب�C��I�[XO"JV�T%���.���ēH蜲%�څ��T�7���xJA����s�������?:@���z1��<<>�S/�0�v��I0trVT*H�W��\�(�<�OȌ;D��iBrf��w`iC�']��ۯW>���H�C�(�N4�P���;�m&L_`{w����ڮ^L��i��M�/�S�����i�fU��Ө��@����z�AM�IS���	�o_�0��Α
�vލ� ��&�oyםLj}��>
��\<��6x���|/���p�'�ҡ\������3��\'�d�4���W5�7�m��(�P�H�Ʌc���[6���r[gc�D��p)8�U@�)XY�Q�ɮe��l���Ӌ��8{�\��� ��ț"ޗ�n1 ��0�ȕ�?ǈ�T¹�����+X�2�(0
����R�ټ51K�R�Z:�A2[`?�2�n\�4��h-$�TSF�l���ґ�ƄJ��U��L��48��+�U|q�US%�iŦx��u���mH�=o����g�H[0�3y���#��?���iB�R�t71���4��� �� e녖�L)�l�e�nr��	�n֥�gk��j��O�������289�$��󵫥~l�KV�dD��L3X�ũtC��=���,Zqkp}���d�:��@��"��?��4?��b���A���ՠ5 ��%��� ����
Ѱ���$}�����UXQ�ֱ4n�~���d��ô�dS����A���0�=d5.���DNq�՞'�L��]��퇞yإ�+:��]6���<tC�cE�LS�<�|+�} n�0If��Uk�KB?��o6*,�*��JFzD�̲?��@�O��Ȗkv�_�����vǘ�vXu67֠�������P�9Q��t$C3a�i�9Mcg�Z�'h�� e��ҍp�JYCT����D.�N��;_	���W�-��b�ZB6�x`/�x/�7#�T�(�A!c���7�)���RK^XH�iu�\��7��0�2��-b�_��/	���h���ꇺˈ�xo��c�H�T:6k��5�|bS������f���NLJ�#�d$���R�s�׹���n^u���PC���s�����F)��^�tڈ��g����!_��2��U�pZ����Rt��x���P��|�2�r�[ԥ�'���φVv�C,��݄-H��q���
إ�^]�T�<&�=�n����0+�18�I��AV��x�Ň1u�u� d$z~�MQ�&�g�d�ecU���➟�.��Y�V�c�q��+�G��"@-��(�xbge�KB�ء����+1:L����IAЌ���/s��+�t�%�Ǝ��N�"��p@淪����� �pMt��rއ�L<��=����m����BK��3"v!����弅��B��=�]Wm�p
�C�E9�R�5�!\V��X,<�!`YS��%��k6����3T �����\��G~����Qa9�͸g�~�V(�vDs ��<b(q��)�s�p���B�Q�k���ߩ��S�'��T:��dю�=� <n[r�|w��ť��2/�M����E�wt�W���1nQG$+�d�ʠ��{����p�k�z������&�l��C+�[j��sAa�kWX�	��/Z"z@JY��=$�Oo���EO����&��ꃳ�a85m��7�%¬�<����Aߎ����1��r��l�>��<n�/�=eď�Y`}e��E/@��;���m -&�=��8�kBj�(0Ģ�����q�%��3i�km݊3���K�\��E�6����RV�?\Q��{������S��㻜�`+䍫h��CNy��Z�FcX
3�޽x�V�h������(8��0q<�ꆈ~�2Z�a(�i.t>��*�q1R��A�dɑ?��]S�hcFQ��o�	��R�X�O���Q��
0G[ l�RJ%-m����=##e6b=|��/�ޙ���m��;h�l�D�8Yg'3GQ�o�$�j��s	Oj̈����o����I�+G8���Q�d=&+k�o�`\���Z�X*Ǒ���2��'��� �諳�Lv�V��N��`YIhgo�r�4�J�NN��͊LU�"@���4S�+���8�(�Z�c��+�����t���	��qٞ��IBf΀�@߿��v��*3\>J�gmi���:��j .����-=�1������s˨���:¾_Fa�b@׃�421ڦ A6�~F°tp&�W;[6VS���A�]�hY�]�-U(��7��� ��Y4{������q�$ߜ$ݩ}t�OG��l�lKu��.�+S�i�7��)�� !�N�r��ڞ�%W.'�]��f(��][������Q�����u�נ�s����I��3�
�k)� 	qQ��3/��Q#�W�Srɳ7����3�;kw�	 �(c�\����xu9Y����0�$N�n�
��U�!��^���]'X&{��+�$cE/n�N<"��.������u��+}\�۱���6�U�yk���UWcY975)G��_���쭔���C�O�\v�G���{A_�x(���_����
�$��*�k��+�vn��m��YYi+�vtP-/��4ddGRB����O�{�	���k\9���5�ݚ�|�6{�������x��`��AI�wx�0�-c��`��ԋ�%�4����c��ܜ�������Щ�1��J��z�ݓ�:8��3c(V���0�~���Z^����<��=:�ŗ�Q.�A���K�5����D��cZY�0#L)�(H%��0g�6���0��$��i�-U���+�;q�'�Ԑ#l{�A�:�_K@f[A�;��4	&��@v�YC����T�U��ȇZN6\R#��z�eZ���M�Z���YW�i@����q��׭'��>�f���!��v4 1�����b�L*�Ҿ�����b�ɣr*M;LF/}�Y|kY�/���2o"x����n?�eM�\�T�;�3�*�oU"����F���ea�1�m�j� f�г���O� �vz�E4�7�sׂNi�SI�5���^4��C�W��7_S�fW�}%����sC)O�l��Qm�[�7.hZ�xL�a��xD���Ñ�fd�ʹ������	�E�Zik'w�.�B�pY5���T��e!��|��r/Ī��x�&�KZ{z��d%r')Z(�4�4��GQymh�bʄ0_S�����F����]A͠�8'���j�Y�#!m������&e��j����u^�؅��y�O�u��a�q�k\�T8�l�"���v�6VY��4m���\�1ϫ&�$*�(���Wo���x�&��	�&�w��D@$*c�4A��-)�M۠�|S���k�h8Aa9�aM���(J��Y\P�0dB- ��ʹ]�y�lAS�uYjYg������A�"���klL�$�,h
-����2��A��+D���Z�_���z�-�_#~���:��+Lz�p��<�*EC��m�g*^3|��׍s��S!����$Js�N�+(K�%���X>,�ee�u�mPSڲR�� ��z�{�]fj�h�g�&�%eDV��W�/�ӎDI1o�z��־����� i
���]�ca�I�<L@
m߸�������1}h9����������"puz�����'����!wW���#?	oDTT
!��B}��$��t�J|�����q�4�/�돮0pSƶɐ��{[.=\*5g���qcR7�pΊN�K�?��9i�x&����������G�P�!0�n�IԦW�-�a�Q8���S�7�jՠ���Wa-��&+�tO'�kQW���YSa���1#�l`�7�M�����p�p�e��9=%���b߅�� 3��m_ڿ�*0��b����yȁ�U�Cj^?�Y��K�6��k����12��L�;����8zU�Gx-�F��@f�e�:�@� v-�]ɦ7�����KCY-I�KGM��Ѵ;z�u}�{�ѷ���o��UTn�������n�y��T��W����9)CGe���a��IRƧ���i��8��y�/x���z�Q�%�S��>N��S	�2w�Ć��Q��<#��`�]�!��p�&3z��dڃsb64��OA��f�D�Y5E��*'G0s�G�c&���3p��ӧ��	�8�\|���5cK����d��Q*.���U �((�G��?�u�Fz2X`\�'�������;�*mO|9[K��{�M��H��˞z��o��;^���	U�-Xl��i�����q�n
����ț�
9eˈ]�&�Q��q�]�w5U��M��<L��.(Y^r~��P���+��հ���N�K݌JB`Yk�lQզ�ZhݖE���t�}�(�%[g
{��ث4�o��w	�~Xw�G��S�ٙ�n�H�p�ėdX�&�͛*玖�X��C�XL<h$�/ڽNF/�ݮ �K�]���jL�S��Q�����մ�� �WB��;���j��G���f�j�ӛ�S񁰅(Q93�B1���M�5�49]�f���1$́�h��26�,��:�B�^�/)P��;��ȑ�t�y�zn)j��@�P#���1�B~�ލ8�P���Hr2��Ȧھ�2��y5��!k��=�^���H� ģ�H?�)�wFM�s��Q�쐎v�1눏�|�gڽmu�r��2�k�h�=4Sg�.�����L�0�l9ky��73J�aW�]TÆգ5S��O�xOEp�[A��P;ie����$�"���9K&\*~)9���踋=���vK�V���c��5x�e�x~p�Y�s�M ���E��yk������ʆ0�g�;�@﯎j��VM�t�V08~��G$�f����Hw2*P)��h � ���;�O0�,��0���W�F�!!	�������(!isz;�#b@����l	�*l�{I���ܿ%n&q�߂`��������Q��8�5��'�#I�%(/�6��V����ݛtd���Àc�$eE�ܬ����'Ҝ�o=��m�x1NΧC�N\�A��~�qA�����q��BѢ��CLg�4d��b���0���	��C����K��C	806s�>����Z���ҽ�e��"X�OC�ۯQUj-���֛*�l������W�	�{����m� ����OT�01�c���s�o�q,*!������!�\������g$��F*w��"�8���7�W'Z%Q
��@�O��x(�H���h�F�6v�L�����w�`��y�\I�9m�B-�<�I��_I����RK������UT���S��y�@����{s���Qx�4�V���<�D�����,�@�6�)j083Ɓ];����p��r���\�=�/}��p~�]G�Z�V�Қ�7sS�u��F�^薔���Wv<���DJ@��߇��c�x1� �I6����6t@��o�G�A[�?��{�y�Y\Ii�J����N�>sY^wJ�U����"�楥Tx�{&�~�W��y�ܽ�����͊���ǯyE��Ѱ�GC蝉pA<��tcd~�L�-ST��ˬV����6��D�����U�i��tzbq�35~���Q�e�X�Oӛ�П�j��͉�_~pnc�W��O��M��*SDg��U@&\��%��l�;cJR5q�iƊ Fh�T��o0�-���iQ�ɵ�ñL�Ѓ���m�teY�`F�.w�Π��d1�?BF@��x�Z�Q�`*���=��Q�n��e�❈i�׻����S��<��J��Wq)#f���dK*q
2~7G �����3���7�L��kڐ�z��Q�55�S���qS1^%|�-)
k���
ĽOl$f�3��,��S�2(�3��o�z�b�]��%�%[���������,}�U)�m���F(�fбW���sƌ���C�SU2(�;����5d�) ]V^1FgD�AC�Վ��v��6}gBN�sar�FM�C�E���3�- 0�^�у{������D�k3;�W:@/o��^Q�߷ �56��&`0��(/�ǅ
��V;�����r ^��#���b����8�$nտ(�������/|1wut�2�ۙ��K;ɕ���J��FE��NMW���q��1������A�B1�<
���҂{�	�)[-(k����.g#}�f�^�CK�U�T�����r?��a,��{�����M�٨?���Wο��/f��)uzq@8x�%޲0�z�N�!:Qi*�%�y=��-�L����q�5���Άŷ��yd8���=�0�#b�������vײw�kvF�rd^p!��m}s3�J�E�M�$A�e�)����1��>���C��)�;������C�>\J���z~r2t�69��F�F��0a�~��Zf�k�u�L�q��G�s$�
lqi�W��Ж\C�:'�ɵ�z�ĈO�c�rwpi�7)�e?�D�s�(�<�~��~8R�v���Y��sѴn "��;����~��+ ~0���T��K4���<~Q�����K:��p����K�l������Gy����.���}��	��%��Ls@T���"ѿ2�${�kFS$�����`���S%�G�Ȼ�X
'�}���>]�?��|sR� 8rƆ:o�Z(ji��n�\���}�厲:v�G��Y`5����F���3�w�,G="}���@��`�j_3.�2�
lK�T!UOj	��K,2a�׋���=y��7�ߝ�Q״�Ԣ�	���I|=P�m;0��^Y�,)�����uFۡ���kŖҙ7�
}�Z0#$����z���������Ê����B�Q�]���ϳ�1kj��?�2Ճ�*�������\<+*�,<;׍`�l�h
V���^6�Z�BIo�
,�/uz�ys9����E@)p��BT�3��h��-�OOy����+��T��(��Cϯ��p�}���V}?����y�S�խ�	3jɣ&4�Y�~ض�N���v�W&E]zE�\Bm��5j��#���Hm�{_��O��S�{��IXW��gEY��2QKE���u�^s����t)�i�~�[oN-��2�!G�'�B��Y����E]ש�TD̖(����(���Uda���I��J��5�� Qɹ��

zT��	RX��~�]�� ��\�ju��ě��Af���;,�M�,��]��< IK2�R_�:��l8��9��7	�"L���uD�|��Y�D3*�*_�㥶P<~[Ď�/'e�k�l��+W���i�0i�Dq��[�c�.Ԩ�ׅ*H/��_�cRW�����	�%U]��c0n-���"�V(�6�FK����"�����^F*��-�ꑇ�UT�c��n?��l'
��5x�V�M�[�����c&#�5B$u��M���s�8�ݩ���ĚZ �j��5u\f�m�*̲�v��&\�>h){A*��Ͱ)$�T�*�P�:��P�o�.�L���\l�	f��M�$����Fq6������C����X~)|mX��6�.ŗxӏ�]��4ﭠ:��]�N0 wYC��[gqP'����-͂hy"D��Ͱ�p����kY1�nI��u(_�M,S�=�{�'7I�W�l�0B����x��2T9e�lC�8�hG���j�u�C���]�P��	Kp'�IO���\}�jI�)��N��b���EϠ��ˣ�2M�baotR�`�u�is�"�/̱L_��_�צQ��i���)��W���şmi.@��K2��e�G
M@RM
m�ea�g��o�l�.���\�Ŧ����U��N��q$_9?���;���w�4�O!��g�)s��k�� ���k�<Q��YX���K��\oQ�KvB����$�)^(]��1P�W��(�.@�oМ7s�>�_	�Ӱ��������N�}��s������P���k>�����7��W���A�x��5P���^g�6%�3;���D������_�\�W���U�&:w��e�'��wI:!g$\W�K�P�`$%M1g��e�Bۤ�-6��@�Mr;�T��d}]��.��F�ӭ�2�;d���xTR�U�ux捳������q[��ӝG\�$�Gr�G�5��*jD#Qγ4����%D���e��k�O���?Ŗ3��w�[`D����-��x��D��/�)� n�����dU߬=t�ؖ��	D��ŧ�6y���<�R.�.O��n�4��R<L"s��6��9e������(L��ԫU2���_���B.Ө�<�+"a��YV��vƮ�$7C��:�������D����m��Ɜ�@]��{�#^l����D��y'�r⧱���_	T�i�͆��0W
�����q9���'0;c\P-�\�z93����W�>�[���3M1�#,ߛ�Ϻm�%e�^E&���Zdesy9LI���H��Y��@�u�
��	z���Qv\�o�`Lvy��� ��f֓h�(4s����Nn�W��TX������Ző��Ԣh�vVr�
�'�^���l/ʁ��፬J���[N�LQh#������U|�圐�o4q ��al;�+c�d�����Mֶ��vL�	��1U�|�U�@�QĀ)�-�*1�G���̠����eE�����̥�9��)�&��Q��/��j#�@$ߛ� �x}D4w�מ�Y�R	s3ݥ����<���u�>aN�B��%�Ab��dr� 'sc����7�f�=�r���m&�WqA��	�ui4kЛ�Da��Wo�������<ˎ�Tu��t,E��78�&d��2_����c�P>�l����GR�SV~����dNx�Q�����?��[���k�bxK��Q���jP��x2_Mk��Г:�N�hG���oK"}q7�l/�RB�?��mVs�[�:x���Ě6�}�C�-��@� /8\^k���k��#(�Dx�S��#KL��Z����ě�Ϥ�6 �jO�ɥ��'\�3xP@�n:�}��'�W����V_`$��0��x����ټ�(�A���n����΍e>Y���$M�{o$YD�1(�0޹�l��k\�}G�, ��z�����m�V|�xy�>��٢�
Wt���ك��4K�4@Oo/ߜ���s?:�d�������B����+�� ����^��q�b��׽O�h�Ik'�{fq�J�.�tAm����A�3n���ǔ���L��.�ZY�e C(#�@����)��	D$=Dn)fm�"����ٌ�Z#-؋'��&22��DP0�byM�CI��g��V�y탲_��d(����>���5�j�ޮOs�Nf�>���+A�w����O�r�����v-�J��& M�fj����)+߹��q/2�[At�ƹ��q���VR���m� �N�Ǽ�[�'��Q�:��U}��j��ki�����F��EeϩF���������5�w]v)Cl
j11�#,mL�9��$��pj��q��aH��3��W��9@t��]����We�¦�	�>ZhD�Rv��Q�o:U�s�e�v�"��"{�>7	��+����D>s�ң��F��EO�U���%w��Zo�5.����q�wβ�-�>Y~�C+IS�:!;��k�9?D�җ��J@^��k�z�j9���MR��7O)-KUU쀯*��b�I��C�
���qɹV�o`h�@�k��s��K\9��4�X�+��o�*� ��L3	Y \̑d抦������A���{��?�_��_��+�-��%����.��廸4i��üQ&����PD �/�%z�_�]�Ȋ��3"���hj�C�}��*ګj�r�*AsH�I���[�0f�G� ��|cۇ&�F�J���߉� ��AoP튢E���N�]�	w�+�������ZH.��NRZ�#��淔x5�9f���R��;�I�G���Q@����S���H�wx�������q%�#9%�g-�KʈBv �nq���hӋr���?�k��I����2�h b=4F����Ab�H���ٓ���А{U�!���a�}���@z��x5ʮ)r1Q�rj�2M)�9\�����u�Y�o�Y�����'�pLJ�f�w��3 �uJh!r�ʆO����~΀��Ǻ%��!�iH��nmd�����F�oV�C�Z|�`�uQM�E�z&dL�ܛ�,2���u<<��Yũ�%vq��K5:&spS=Xe��/���M��i�$�E�J��J�&Z�O�x��J �̆��M���N��i}FԈ�-zof�4������Mۤ�-��OK����|=!��q��E�Y�MPL���`eU��u�����	`���שu�\+����f�ɽW
��HO�E������:<^vJe�e��k�M����(n����.x/>�s���m��q���/Gχ���
�K6�7��6�I���
�rt���~|Y��GJT�����Ԫ��D�ê��I0�:l:(l�'Ѣ��#PS*R���H��x���m@�|  RE\���@A(	��ʔ���mdA"ο7(�ճ�$g���^�Y���k~ �������n�`�!o!8��n�.4"�͙�b�W���8�l��؍N"9J�Xe*=܎Լ��	~��r�_vs��}cn|��Ww�_��%�9��:-�3��k:"�1V��(�_]S���3P9=��IWd�%�H������$S�&ox���t~y��w��|��<�ߨʻ�Mp�����;�VLE�h��v��(zò���aܷa�"�} �v���%�"ǎ�iMz�*������I����;gG�����/�JI�׸�`#6v7�2w��Q��h�����Rc�p���*���3�a߫���9��|�rv�>[���$��y:`�B�  @������6���л��Y5���t���I��������X��ͻ޽ju�}�I�h�q0��"��qdl8��4|�-�W�$�r����Ն�eRUlW�BN��>�v��3PB!s��)�:�����P���i�~8z9�ĝ�z�M-���G��{.�O������JU����ݾ;�#ynL%����Lޯ���xX
���N3���.�����mms�`/#,K���2=���{6I���ԋG�\ͨ�
��c恎����*zY8]��˸��y��e��l�7�[Cd�����6m��w�iS^��g��>b�cc	|j�RtA�#��0�!�Ô^�l�/'�uC��Q��M����Y��W���%��u���17O+o��v��:�G��H`u��1ߝ��ǵ������v�م|�1��@�����v�Jy�a��"�p4�\7�D}�tXAnR��(� �U4H�C�v	���_߮JS=�N(�a*�S��A�W�V��M L�t�����3']o��z/�`e�"E}�^�t�u��o��4�8ᏹY�a��+}� l�3�Z���V��n��U�P�g[�{�� ��#��U~�6�
��N@3�^����m��/�n�?Q*��d�.$�^�~>%w!�c����`���\�q:�3���7�/1���@��~��_{�]���Z��������=���0��e�=�W��1�W=T �{V�+�lܤ @v���<��$��p�Y��z�A�yZ��
�[3�����N)���$A_�����H�\�Ϙ��%Γ�{=l�U��´�� v���x7
�F�Pwc4��!�$,-Yoߪ8z'�W��*�:���l�����E��gz�"��X���xmNJX�L�����$n�q�J-��xb�=����6U���wD�@�B=��5H�Y�k�֦^���������2�c��۾��;�&MiI��T�vZ�HH�ix-��ґ�w����?��$���gϪ��Ǔ��p�D���O'�����Y��d������ʛ��} ��j�)â��e{XA]Z*�$�A܁E��:I��)��|���2�����xsle�h�Ǔ�IJ����>���f�JH�:��H�䏆������R�g�_j�2�nְ_r��ЄK���5b�Ƨ� [#��@n�T��d��7�l5���GV��aթ�=��,ǵ���BV�AS�t���@5�?��zu#@���~����_;j7��쌞%�s<8q��c��x�&��y��VnZw�!���	{!}ַ@O���&8r��Q�kC�;�P��؅����=WId�P�8����[5d'ߒ ��ΧQ;�;g�"���K�7@p�ad���)����2�L�5e��������hR�?J��l��K��w�;��_9x#�2j
�c��������@���b��7v�E�P���[O�5���aވ%���#�Ɗ��^���7y@��D�M�0	�;�}����26�m�)�S���6��*,\�A���.��Y=(*FI�밻c����x�����
CAŨ
^p�x��Ј1��m�Ak��A��U博Z����Զh�9�D{�怇��tGS���\��#gLFY�Ɵ��nQo+�#�#L���]1葽k�Y����e���r&�"$e�A���I������䔺W�Ȁ����\�S�!��f��`�I��tY�h�(|�j��<i���p�{e�o��:bj�3�͡�ZnW=sk|�822)��5�vz��f�H�k����� "��`jAb�3�`n��z�Kq�����������5
����AM����qj���)�s�WV!��*mw�b� �7�r`4�R�L.n�%���P���)��G�G�L�䃹���� �[�M߰ J�����@�C�X�,am���M�?�R�xt��3x�q�[S�V)������H���Ds���m)�/��D������ݡ�T�����8�Qǆ{��Q|Ϲ{�ą�Dݮp�`[v�e#�P�k��xI>�Q	�9�@J�|�	KB��(��}�t�w�2e��9k�U�����E���kz�4�������*-�%�U�*ʱ ���I>��7���������d�%h^ܺ9Yb�.�fre���X;�. ��7��7������;�_�ތ��4I6����k�2��]_��GV����*�i���6���}/b�
>yv��������'���k���*��$��!�����e�!�1�?��G���o���f_���Fɼ�/+���gy8�A���9��t.9�v�*8%�|MZz��>���i�Xo'Y�b!��5	W�gi���	�1z��q8A�M�0�95ߔ�.F���!�@è������JZ��P��LX�~暘�u�z-�U!��K9~�n�.��Ԉe	�|��r��-���0��15l8{)�!65�߽��ڑ�Zϫ�o�e���!4��%�J�'�v�l :�as����id�L�q��FNҰ�����2!�Ȉ:�1��w?XPT�'�ߎ���v��L��[MM�T�ҌA�B�;R�5A�h�d�񖧸����U��c6b��fz0� �Vo�����Y4�:>]�&FM�Ⴠ��+�:#���� �0'�A#uK֥䷳����NH^��/�1��t��%}tQ�-^��i�-���!���	Gn{���%4�y�`�Ր}�U�T�#@�x\�b?Xy7�w�R��o�;�
���{Ak�x8�� O+M�層x�*hΠ�U^�Z�ɵ+�Ԣ:��q�.&�
��p��6��H o@F�F�d}n��7��!ׄ����$���$�}2�Oi'�p�󻧭����%L�X�n�͂A��϶S`�*�G&�`�,��%g#>�
Y��l������BR+���H��J�\4YDҳ��v���l�#*��3~TU,��@ժ�������c(�Z��Q;�(���T��R��y`c�B���3�� �OXZ9F�yJ�1��l���/^��Уm�@y�/�-�²Rq�%x�i���QQ�s˶9����N�h���՚2X~y���'\0=IL�gbX2v��+�J�����_������Y��T��W�LO��ы��nt�3@sĠp��X�+~|)�c1���`�tz�����X(��j2�d�*�3�m�%wE�B�D�~���WM��
�w�IX���ӕ�'�r���)\I�� ��ڠg�,z�F,,W��5�
��,x��e3���N$��&E|�h����~�d%���$�?��{(�F?��NӇ�s
z쒇�E�G��f5��X�2v)���e�
Ĕ� ����swt�ЖB	��22��h�y%߁W]?��e����~�#�����S�+23��Ȧ���!�@���g)��L�h-7@͂���6�z;�UH�*ԥCn��c�?��q$���J�,$t�:���I}x^�Ŧ�h����u��O�!��'u
?�����ߍ���]ē1#���Q�\/(\��}��4�:{x�:l�9A�����>oEH�L4[�c�kk���/S�=�&␲v�.��~|4þ��U�!�.�^�����΀�36�od��a��R�Პ8r8rO0GO,���7Sa�����[L���GW�y-W�' �I��,�2
��6ܔ�g}��v�w�s$piS9��Ϗ���J$q&��I������_�媀~[�Ǝ�Z��A��3����!�b��>��ɞ����O;��8IL���ګʲ���;���j;�go���C�Ǘ��T��y�ሶ���Y�{��
�G�H��aLm˴�vz��5�w΂��H��Z�@?,����t�s-q�e��l[)�h �B�;�?S6Y�����ex��,4����-p$�I4�rcFԴs������1'!4�E��@��Q��>M�!nOVb�%= /����L���2�^��������Rs��c8\���R�)�!��hk��0)ZQ
�rڍ� �^�`�ri��#��ؚVԬWr�UV)������Aה~�4���}�oP̘P���}шNln���%�Z�P��t��s�<�Z�wN8*�����q��60v�aB����|�ʒ�(u�HWTK��=�?��~f�`Ơ)���ާ��ԭZ���yy�� ^/��m~�i9��
x�\��P�Ǖ��[Q�9qc�%�HJ����?��W�T��������IF����*�,E��_��l�c���U!�ӵ#��i�`�k�.q�8�LO�5}�&�H������!��AB|.y���b��,i��m��@���� �ԣ^��
5F��Ar�Щ~e����s�v[�U(�_�!n�wt��;$b���G�c�V���Sa	��}��M���M:�6�"�\<}�}v�J�Q�rI". G���&͘x�ZFb�����E]��5)97�������^Z{��9>�}�����I�q7���lT��Ա�H�Ħ�qr����ié"ʈ/�N���t>�C�;�alTS�s˅P�J>&����t}16Z��v@(�j�[k�7�����)&�o�Ԛy�(�3J6j��].�8i<����012���Rk6~����\��+!���dk ף���c{Nu)�=�� �	���:�b��2�0�\�М���?�Ox	�Š
�j�!s���=uܠo�%A�	|��D�׻�3�`^v����EW+��[7����=�;�ox���+x#I���+�nw�K'�eYYƝ���X�&���J���=�&�V뫭�ͧ�/�"��7��*7��6�>v�$��(�����R�@��K�Qa�早��+�A�W���`7?s�v�.L+ytfӲ�x|uIo�2���]Q�\O$M�cn���濅��ӳ���(��T҈��kez(��\TvF��X
��	!�T�-��՛�#@�9��j���dULw؄���* #!��P��2��V��B�-��K(�����
�v�X����<Jc"m��_X��!���%�NR�k��dm� )L%��ك�W���}9���"��z�|�A���Eb���e��D;��Fg�V�YU+�0�$��#��՞��H#-�`z�[���<��������o���\y�w֧��6�������l`�g�C쬼f�8����Y���fMˎo�.j��Y�wSto3ͅl���-۩��9���!�ԣ�NA'�Hق9�R�ͩ4����M����M�j���� \�P�i]<^8���^�����,��0%lB+_g�#sVq	-��{ʧC����0�d�O!d�u�СLÊ��7�wy꣗�=zV뚲����x�(G��I�$F�99/�oȥ�4�[qx�%E�~�=h�l-�!0���r3�.`��XsBX�=u��x]���e�a{]0	��E]A9s�l|�[��Ʒ��m�_�v]ZK���M,.r	z��W,w��똉NT{�(d�BsrG�S�~M�h|��9�Z����������鰃�F�F�g��-'x��y��X@W7���g[ٖ�:s�|�K�L��#�5eAo���1FA��T�����;�5��7���j%u�W�8�=\C
��!�jEe�f��l/�RE��;v�2�OE����h9]GҬY�-�P���)^�b|�a)ƬKG��Q��h+ϛV�������T��m�j�<'��xhI��`�#{$ro���(��07�Q=ڼ�8��	�4 ��@��A3��v�E�j\��2��b�8/ldU����&;F�I�ݟG�x�9�zt�?��p�QQ�,��hM^�=kɴ�P�ZC���k���i�gs'�r(d����Xea|��l�1�Y18��36�����ƒ��fD�*�ɟ3� )���5�F+:��>��B��O�f�٥�J�SIa���m#�e������PQiP=͝J�"�u�t#w3��cyA6i�q�
��Q�;Z;�:�U*#zO=�8v4�`jU����/��{�o�_ �	RŅsre�B&�~�<98���*O����ǥ�S��t�v̸��u	o���qŞ�
�֞��+��*��`��P��?���t����Y�#�/�I����R��$^7����|c��3�N��Z�称�OfF$)&���t8�~ⶁ��EN�#��5��Ʒ�DBF���.��7�'��n`��2�z0�ڃ1���BXq PI�ΰ�ٳ!��q� �� V�����T�C׺�y��
H�l���6�J�y�����_S1���|��
`Z�� Y���WH�L���yT1|�f���T�N�]��%)r���\H�3DoK�<����a8�)>#;��L>M�b�Nh��E����Y4$%j�GR�R;5�n3���z��`"��I_�+�"����6�_2���f���҆��5u@���~�4L�j��:J�+b,ma�q۲i&1�H��s*���ߠ�����)z��b ,<��K\���+�C|H��d��fRZc�	��C��X���b�$ �YS�W��ir�JV��aF��|�t��K8Z�̜}��������X��w���N�H�աK�aR�DUT~���|;�$b���P���u��O�]��H1(#Q��(}bh��Q��d��ZW�h�ҕ�\��D�2��$@��%��=������Q�G�rB�s�
A_H,�����G%���>���6il쵵M�J���l�ć����++�(�aՂ�Ue��97�����bH+����wO
�`p���w�;�$��Ҝ��JX,��z��`��b1(��x*=�c��)|;$e4w���Cf}۬��E�2�nC�X���\"fd��v1��O>���;�[ 6:�� ^"���$3NRۙ�4NB�O�����'���Q�{P��V<����?�r�O���Ձ<����4<c���V�^X�GB�̚�O��0���TA�z|LZ"h8\��Tԕ��Ə4��l��B��an� ٽ�g=�N*8�7_��s���R�V�ya��-��6�Q��*?��7��0w�m��>L�{��"���?���v��L�����b�-�����=�����>"��RY�y
Yn@��\(�>�KR���Y��҄���T|J��X:�U�Q:CgɸPn�@��.r���$���8�ec�qd�����D��o�p*R\�����2P��ϖx���լt�'ŏ�3v�(><	��a�z�"��qA�?B˯��圵kl���z��Nq�l�*�{1��k6�D��D���"UDNݾ��ܝ;u<�a[&yj�m��������Ñ)�9ܠO����OO��g
]��G�̇ U�������j��3�������>$�$��)�:͹g��H�r*�zB˅�{s��t���bL��H�����Q�;�`=/��E����E��i�p���Y�]:�a�ˎ+P�Bm���]�;��y'�V�Wo��;@7gQ��9�9<�?�7ێpd*�&G��;��ԭ<r¯����Ѳ���OF�R���pk��;� '�ʹa{m��]P��0 P-����XP�ReI_��)mֳ�V׀Il;�����@<5��7Z�,iUW�:��-�Ŝ����gN��5��ѳ|8Um}>k7�G��Z���@�2s���]i�KB쯮�j�5�����Va̷+oX�i�w��1V�ݪU�%����\�
�KN2	���ev���R�s0�.������<c؎T�g-�� �]�4n=.%o��B� ��೯���ltwk����K���+~gH�Sۅ%�?�'�0�ILˆ�T|dȻ8�Ϯ��H�i��?�}�g��DHYh�,_]Sg*Gt N?��KDA��Y)�<⍕h���i�壘C����A&�(b9�9.i5�l���w�Kҫ8*Y�PCh���j���j�u��@m?�k�k�ٜM�u�e��3��n�M0��r�R��/z�����I9�/��.k㫙�/Y�����ۋ)��u�t������DI�Y� ���P'��d���XK+�r�i��f߳�����/�pHQ��1fW(;8 ��d���T迁�*��V��q��'4��K���B��|���ٚJ��0���2��)����w�-��h�P���|	�3W�w�Yɤ�^��rNp�SZ�抩I�e��6ܒ���;m�')����2�(�ҫ�,�����M,*!L��#!���Ȭ�"�vd��Gcu��B�0;��� c�(�܋? ���1d-G�߸P���!�Z�Kq��M���2p��}�9����F�܀�s��|�����Į?1Ȱ��%�ֽB��
�y�?�7�c���O�-���d��|.ﾼeT�;ۯ5nq��|c�4�������c�o��y�(:PU���Y20f������� ���H�=y�Yn��{��^��4�j 9��]�R�L�ExH^I�[y(6�:G�n���������Nظ��ʆ���mY��!)c�uPTw�	f�.rN]���o���{Fi�}#^#o� l�俷�x�s_���.�j�o�����2A�ƞ)��)��MU� q�4'��� �l���׫����9��!n[�S8a�)�2^�[�%�^�&�D\[�@�y��)��CZ�����>�������N`慝�n���v���Y�̗�W̩����y�k��kt������|V��7P9�]$�q�f�Zk}4y�j�1FrU���h�7��u�]G�m�����S-�:T������������/��N������6�ӷ�o�;tKš�8'!���& �,�2;1���ْ�Rj�|��|n.�_>^E%J�e{�?:O�$��o�lW��P�u�4V�Dܨ��H{)F�̵���켅kGu���B�v͸^!���#����>�Ƽ�C���c��
c3YFW��2���� j�O�*��*�TI Ͷ���X݈V�b���U>�sg�+��WY��ٮ�;�ɟ�o��Xq�L'!l���RﳷX�G�l���*"bϗ���&�YyT��`$1�5���{��cc"���SnW�"| ���7eqe��pV�W��j�
t�5B%�U��Ǭ"�D������{vt &��O�H!�Zd!|�͈�8�=�E_�2�h@^�3ɩEE~�\��W��U��S9H;�7��drc"٠����ؼ24X�(���C�?Eː�S���}}�!�1f�2��?�Ue!<?�=dD��лq|i�=��l^��v�������.�#��X~!1+P"���ԕ���K��G�>%J;(�@ii����ތ��Ǫ��~F�}(B5ȁ�.�6!�->�O
�:��>�5���2c	Q��>��0��u��7i����\�-�բ�:6�žT�.~w
����6�-��c��b����ϑ�:�!����C~c�����W��,Б'��U3!@���YNZ�����_�[�3�ӎ�=U�'*՞�q�Jy�/Mr�}�F6�iI�W�=; �i(!��j��7f>������ځ��O��jG��Mn=��]���O͛��Bp������C��|��3�DX�%��������<b�x5cu�7�]0���F۵�9'2��;]�"���E��]�#��ȃ��{w����t���T��H)��s3%�/"��� s����4ѵ���/Q�)E�I���%ʳ;�'�z�n�j���s狡
����(h��u ���`��"��_r F��e�m�)w�7�؞5���^"[��s�&��I�f�W�̼s��^�ۀGp/ڲ+�˾��(:�:�;<cx��O���,Y�:��0�p�喡.7AH��\/~e]}����{������
FGK�����YXF=�N��Dғ���Ht���|�� ���I�K�|��N�J��� #ֳX?��ܝ����{�(�pdW�)�)���%��77����O�[��@??Sw�EC���*	)�>�3�����kdT����
o�Qq(�)�^�ۘ�Q`���,'�G����O�V��v���xED�@ %�l�H
��SW-��}�U�w�U|<X|�#��cZ�����#�'vF9�%
��I��V#	l�^�:�s�\k�����c��=�bB�f簋�`�������+�5d���$\���9����/�u�B={iE�k��*R������''GcC�N�4��n�D�&䡪]})���`z����;9|�u�x����m�KͶ��uxc�~0A+�	��6�����3���e�M�T�����#��E��"9w�����!SDM�� ��Uц6����hB�P@T�?����)z�x�Y�����j�H���˂�d\/�PV�;'��Ճ���PG4��NU��Z*�^.۽v��l|�+�<3ˁR%@�>����(�E�$9B� �߁���m2F�l�Qu�d4��Zyv��
	"�D�s5|Uq��+�f���؀�+
���<�N��s6��ܧ&<�;$��{�H��[Kjny��0��X�뗖M��dk|V��G� ��Z�2�Al����I>�� �~.esd(��Q�����;��]�H�Tn���|�.�ѡt.�E$1�z�2���A+��z��>*��̺J,�A#Y6a�#�+sULp_����b`E�{�� ]�"p̅��s|����gx��ֈ�q��|���p�T��<:�s���%
Pc�5��n��8��4�_�M�m�}R�o��n=������� ���e]le�����fAש�hG��A~<X��*�6x��2Cn�Ap�Y{����QNHc˃-b�j��t������c�&;��Hv�����a�Vډ�L��w�η���b-�O��|�*OFgG�{F�`W*Ř��!;3�&��(�����n@i&=&; ͸0*õ�ƽ�c�k�`73�A`�����`���xbe�$���k�:VH1�s~LOR���<+(%��x�@��,祪c�L�	ԅ�r#я�	B��0{��q��>A���BQ�j�A����2�Sx�sW�
�r:l@0���lLF/�`%>�����6!T�V}�0��ģ�+�)j�7�2ؽ&Ѷ�4b�"�ś8
�j�Lk�5��y,D��U��nP���6�j�2h�h4�<wx�W�H.t,�F���0Ѭ��@	<�ܡ[�27�f'��R*��&@�<�
�|R�=T��r���~��𑩠����x2�I6;�yM$����q*A|y�>�;}e˔J	3JV���b��'�Q!���)]�M�GL��s� �#tE=�==��;d��oҎ���{v���BU�����-u�F7"�����4�LyF)�к"{�
w�(�u6=Z
������� ���a�������1�aR�WL>h�j��$�_��=J[��q�܄͚d����0�Ჶ΄D��Q�����A^��@���&�uCC���_�)K�pִ	���4U���Ή��U�L��F#{<Ĉ�F�y�]��Zr�[N���6C� 4G�Nx>A {��'_� �w�_ N�U��y����v/��4�����o�	�'�ˊ_(�*$�?Jm�3�e��$y�c���:.��(}:���ː�i��]ԡ���bw|U A��<��
��7c��Pv/��m�W�6�)�j��J9�����!f���$�W�»����xLB�c��+@���6=<�F^R	�5�?Y�:���}b{b�%Tr��C�٬	���-���!2e���z�M��g����kZS����������'���)�o�/7�S��l��70��4�\�
�V��y9/��#�g4������9�:�5n	����dƟ�
�{mYA����pTS�ym�?���h�P�.8p�����paK��E�4Ʀl�"v�]0�l��*����0�<����Z��-�.4�����������X�M�y�$��H6��4C��#ۜ�C�D��׈0��"�T���'��h��{�l'�*� j�#9�:��0`��*��U�������%���a7앤�<�O��"9(�{j��kp$c�B�͎ks�:CJb`Q��@��ua7'M��'D �#,G����3�%����(�G�w-���m��z���2�Gc>�[�E5����e�i�mTh{��m^�U�L&?1�E���L˧W�9��^��� ���j��z�A�p*|�}x�
�ݓv�D`�OY���{{��t;��o *�e7�ƅ$C|W�;�T�g\�����؛b �����e���_�;�k�A(�L	�^�5�S��`~"�J��~�Yt��kVt��˝��Fp�]��e�h=y}s$���u
!�I����9�>�*m5�̞<לe�՞�}��H(gp�u#{,~��M��2 }�m�릷�b�~�w��'���������R��F%�Mb�b��>;3�G���lC~	^M!<�����1�{�
�}W.�[�ϩ��7�J������GQy�k≞��@Z���@�ȩ�DA�a$�\�!6?y���V��K+���)lSvf�?��'��c���~J7Uy�!�20��}�<G�E6s^�ߑ 3ԭ��QT���^�>#t�b��H����Q�Xj���+������D���B�_�x9��X/�a�ӡY�	{L~���;6�>@�������,����L�~��m�T�3�x�qC�uo �1�z�����A���mDy7mE�E�p  h_���k)�	�f���8�g7��A?n�F)bV��Dk׊P��,�~�z�d1����Ӛ�z2n��|���j�V!�u���6�td����hR�_t�SԿ�0�㘻��T�WX���K�/�H�uiJ��:aXȠ��L��gٝAq 9�����^��5����B���؈����VC�Z�I�zU��|�.���3-�O���N�����px��͎�~�Mu�~� R7i  e@�8���<s�cdt�HYJ�$�NPZ����[�����rX��
�I{�]��0�9q�k��.���j�o�P�O���F�;��Y1}����&Ҥ�Bbõ�%���z�?G��=��G ��>=���N�Zs�{L����/��@�L�ܓ�]9x�3��Z��;�����m�n�.P,AL�Ҿ���/�X^� ����dLO|F
A ��6}���p_�������G����H|�<���,Эiλ�r�:�!^h�J:V�����^����|�|��������������^o���2��B�n���sOدff�)�I�%������n
��V�Yy\4
e�e��
˪1�QC�=�A ��՗��F�x�X�)��Dm�c�k%~�.��W`����P{ ����I/ȣ^/��W6�fL���Ǣ���;��x�3W��G�N�N����xT�P�F��3?�j����*Y�Y�W[/��X|4Jɫ�����{��v���H�%@>��;�]��s׉�����^K"�upCn�}����eGհi�?.�@d:y=o@���R|�m���,����P�T�2ؒjͻ
�)���6�G��E��sʦB�R�0^��}�Z4aV�<N�}p��Et�� ���p�/Zg��'հ�g^k�y����	��r�7�*�3��<
g�* �"?�
�_A�S����Gd�k� �>�b ��A�3'J0��O�>]��h�ׅ߃��ChvE�5L��ƭ���3�#�G��M`��&�S�� \���aʮ�9�y�̕!�cu�5�S��C���u�F��qM
;tB41�w!iI	�2s�IniY�.g��;\��d	a68ޖV,4��$D>N8,�*�����h�[t��9�ڭ���XWС0���F��P)JU��:�����ܼ�B��BEa�_+%��`b#jn�-��e�7���}��p�F�^�{�����L��u3���!\��R2{�D��`]�:»	ļ�T��5�0��7�Ty��.���<��t��:�ќ�R>x����u��7�9���6����{\�b �l�φ�B�yϊE��!�]��f*���ZU��H�\Q��S{-��3����M���P���7^G��I����Cܮu�</���:�!S�x�L�
G���iU�T
��=ʄ7�i�Gs��۱����l��$,��l(2�JW'�l�c�<8���8��-�vw��x�������?K�-���ֵ���Ϝd�.���C�T�fk�~cP&u0��B�\���E�Ѭ{_}�[�h��q@��ƙSV�.Έ��3P֤So ��̄�Ҥ�|b�U�j ��%��o�	��C�;4�Pзi�Csu.<��Ze�C�2��E���}kM�Ⱥ�rM%=;�v�HB��p;=�x�*�@k�]HMȻ���3�p.G�9�l�8QD�T��)�_C@�w-��a�9�r�7�����Og�VM���tٸ3���:]�b. �)}���=���ɗ
�ˢ�[�YbwH�Zi��|�b�rC�eQ�Y���Wؚ�a�P��z�*�Z�� �1��J�d�áY��۔i��r��p�nb$Ed����h��SU���[o[$��[�����nD)C�!<�FB��`��z���RQ��ݶ��4���N gg0\�#����>+m��,ic[���[h�Di5��>L/=_��$���`	#��7�M�6��U,�<K ��#�9�9RZj��!�J���̵����Q����Zgt�[HEO�HrI��,ܥ̢���P�(��^����h�B�*�L�\P����x���H��د�T�<5��b`�P�V3�7UւD�;�"ǭ:@��cM�Ɗ2V�t�G�gp�Z���{)�-ϩ���Q��B�0���U�n���!�i��4���/�$]��v��a��.��]׈��#8ʁ�9���d������r�8�`� ��ư����갩 �{�\$�������ffu�Ba��Bfx�����LR�9��A�_�z������kХ(F�P�����Z%?Z���\X�u��s�x��9�/ژӳ��ӣ	.K�7�ED���dp���خo	c������G��80ZXe����z���VL���\�������{#A�#�. H�'�q���k�	1�����(��ߛ���L�d8jq��a��:�ƒk�]nm�g���j?��R�(����?��ʄ/����B<�4����s"����pmMt��:a�Y�1UX���;�Eᣄ�)%:��cZ�M�0BHt��0h-X5�t��ws����O��|/Cu��{"�k�J/��^Δ�a�{��[n`�Њ���M��d%[Ye��	47�V&±A�43%pM=�N�>z�:eKf �ךy�J��G��'���h��[<U�v�(�E_�:�`X��][�}�r��v�r�~`c�	jI�1'��bV�$�"����n0Ȧ���&=izcn������@8c��^ٍ�����F}�{��*��R�I~qk�\��W������ώ�4ÃH_��T��t��で���l���&ק��&��pr���պ>�!��-�d�x[)��c�d�s�lX��~����c�X�e�Nj�8�+][��������ɀJ�!� ��6��U�y���Ys��k3����P��n�/�l�$ꆜ9?�B��J����s��޲M�\�ڒ�&��]�g�=A΃��Ri���6�~�6�|Zs ��A���C�Ucgf}�I��E����}Ú��̎�'���xk4�F�DR�:o�=1j��`v�m��t��+����-���wq	^�d�ZX~d�TN�P��LˬSw����D����>��A��a�1z'���O��[��L:7���	Ig�#IB�R2I-��_	���hb 's��s�2�������8 [��}Y%�Ļ�zD7#@O�#�)\�aB�>��7$�^��4��Y�
Ԇ�T��I`k��<�.��gϬ�P����ǝ�v>3!�M�R

��4�H/z�8��Q[����7��h�Z��z����F�,�E���In���`pJ�*&GB�n���پ�^��Zčy�q��|ɣ$�W�@�@����G��gO�b� ��nuO�А����G�&۷��}+���P>�����	1��:��J}�ɵJ�8���R�:)a��ߚ�H��B]P �&�0}�
���R���$`<sZP{�Z�}�[���T1%=T�H�Wʏ9 ���Im��,XG�x����y���S^�y���P6���y��Ī��B�c����+�q�b���y�(HX�"/{�{E�Uu�O��p&<�p��T�j[Η�m����<�$R���:k4u�
�<<�8�|��,���6d?併ݸ-|�VG��JV�<�טBZó��Y��MԒ�wd���ǈ!=��?]�^ ��[�3�I�K��G��
�,Μ5�::���e�/��le�u�C
D��8A�Mr��V���`-�DG�,_I!m�ZqWmI�r ���,�!5:��SUm'����6FA%9c�($�,/-d0(ٍke���ݜ�n\a@�d\��L�~��C7(>ej��̂��ʵN}�*�wUHE���ґ�O�=�X�@uQT��3�s��=�o��k��&]uLl��!�`��O����	c��A%��ɰA���Ƈz^�S�'v��Tv���u�\=6�V�b g~Cm7ɛP̗�R��Á��$,aOT�)�ެ��|���hn��|l7je��mz�/�b���ie�F� ����bGQ��MmD(10P��Q	�� �f�Zrj��hBYp.m�� ,gV{4��֔ �&�y�}Z��� ��y6��,YS���g�'��"8{0:#)3��tc�n!�(�^T��A�.1/SqϷ��J�#�~Q3s�s����@��N��ҏD8��,����_����2��m�~C��D�!��c�~��S���m�7�*�@��-c��;z�r������_�)�ɛ�n�3 `7���B��5��Q�A�N�a�;�L:��'���O��|/<*Š�������ތ;�����!_Af����A������\F��N�('`����Ͽ�}/X���|�風���<$�t��i��4�t����i�� 3�|J�F��x��C��1�CI�{�g�F2k�U�|��ki��[%#���~:	�Ҷ���9�~��TM���0I�#
r�O�o�"���M����\Qژ���{�%qċ�*�uH@���Z��3�n�?j�<O@!���j1{+����TROyg�3��y3K������c�L�u�Bc�5D��#y5Y"��ZN���7�Z_��!�?����6w�;w�wg��&��#뽟�B�=�A	�J[	�7cۨ��"h���!(&b� ����_�����p�&�q��]�s�"�z��E8��7�9w��%� A����_}6�3>�D7���Z�7E��:I�Mv=xK�Ŭ�Ir	 ���\@cT�f�xވu/�Ҵ�R)���9/��aڻ�6�B�HW7֣s��<�H����EN��7z{DQ]'H0���k�Ǳ/N)"�����,�Y�jXXuC��1�AH�4�[�U��ʁx�CD��y/v��S��/���H����e+}�7��\�(��T|����-��}v���#�=*�W�y��������4R2 �&z	~h$Oٶ%��7޲G�/�BI��|"`��kJW��q��,|n3 �l�����eLܘG�wS�M�u_U��J���kv��l�u[���7E��Wmm���Z��k�4��	� �3O�ZWIR������1Ƅe�L�ݎw���$̈_��E/�ғ��Y��+z��>)�,��R8�Go���?���N7b΁����&.Gk1�"UB�j�����pk�x��S�[����~������V��b�¾4��V��fV�$�c�U9��(!6������ɣ�YMHO7�ܡ���ߡ�Y+)�nc�ʨrS�s���̨���@�v�K�'����.�dr���i�n@���X:�5;<	+נ�}��v �p�De���<E(ip�-ATȃ�[
$�]x1F���̭K<C�'Qڜ�����L>����P���]}�����۶�_a>����Te��Ũ>�}o���%�vʈt`+H���A[EK�9�ke���}��	$�B׌���Em��l/��Z����!���&�~N���<��ð�J�?t�;�t/�����H}g��9���Y1�����,N�ssf�h�(���m����f�����b�eV����C�����#09!�a�*{ڼz��\�'%T�L�i�w~J�;�W�-f�h䚄[�F|��/S�e��8�6�����UX)���k'�]���6e;+%�t[N�������!^�<��G�p��F7A~s)W���R$f�A�Cf�|�&�i�#����XCNRT�P�ܥ2�K	����2�w�����K6��Z�����`�/��l`n����O���@�7ٕ6�P�R�`��U'+_�:�x�7�xhf��,��ud�#h���V�*�̪Ĝk��s�'�j�U���|dX���dY���A��=��(8�-�l�W6Q+DK�C�o�+ǻ�O��Ę�DC�aL1�Rg��f���\�Pwah�IkQƶ���m�z���+E��U3�g4������ -�ڶF�}`�L�Z����BH�Np�5F8�O��b���1�1��uU�Ǿ�eJȫ�R�%�"4Y�ܦ�u�c������w�3�փ���4�#A��mc37��p�]��z��tvq;��.hu��8���,Ғ�S�U������P}ft�=��*KE���^䍝 �ۖ��?=l���f�D�=�r:g��4����o�V��19q�{��R/�Y�0]����`���8-�����������dK���[��yT);����N��4g����6{��F	c��^4T�&@�M��y���F��ЁH�]��U��;�����=�g��vL.�l>��/p�}���,#R�6��	G�Hc��V���U$wO��ck����.1 jDD�(�%��$_O���zl3�Dv�vf�<��"��<�I+� ����?c��-Ts��4
4^�"��T�&Q[~]U��W,S�
��z�3ۃ�������o3C]964�9"�o����h���I6�w���eȐ(��4U��].�R��� �a�KNe�ƕy~��ۚ&^�};�������_�7�&���~�����>�l��,�|@�ET��\��u�l�t��qVcv7:^����"���W$>�:ZAcq|0L����u�	�+d��3,�ݴ����˦��z���櫻К���\�H^�ᱸ1�*V�Ų+�ӎ�q4\|5۔�ҙg_��f�]�k�;����K���Nҗ�����e-C ��ޔB>K���O���5G,Қ�s��VZ'gSb52���-�	���D����ڿ��Y�ف�֠����9���r�|Pr��S\�	k��v,�ՙ�2�H)0���
>w��p�HJI��A�eGm����9�ݴ3��a�P6iX�]�Z�����Γ��81"�7�{�p\q���bdD�U�w��������vM����������܋��*�xs̄��|*pip@h�hҤ�FgqF�|���h����Oؑ^y.���ǐ��{֠����fc>�x(�M�iXcnc2>o����!>�u�'D�b��S)�#����A�3k����Er͐َ΀�ˀ]v~�!��{��*��Q���Us�����+�d~�|���K���Kt�S�0���w�}���YG��C5�L���*�wĉ�_�)<�� �@�� �_m8�s���:�>;Ə$/U0*��ȳ5�����7ӎYp��<���P�;�v��ziX�%P�W'���3�Y����%PYC׸�p� ����-	���7��yu��ɣ�����Y/�A���z.�\�&IXӜY:���Mش�2�R��f"���� ��.a{QT��q����4��Tʿ9͍�󚀜lZ8��-�]��SS�K�t���ُ��V�*ËۼE�3`+KҚ����:S���B#gk�e��z��A�c�3T����IZ$B9� 0��[��C҃�� !��l^��=G�i��Ҽ9����?�;�����5�,����N͇�'	^���o>N��T|,e΍EuP)�I靧��f�N>t����Y����L�r0h)�SD6�V��4�6��
=ϻ�&�OW/�9/��t�T}u-�5Ҹk�����u���ԭ0OՁ�azK���O�*I�;���l�L�������fF�R%�x=HPS,^�݆�J�7�!R$d�!���� u�A�_<^O3�:�q��e�&�TPh�
�*tՌVߒ���|I�� �ǲ������k��'�m��*D8eq��OBT�[�U6wW�N���/��V�__�`T�0���y� �[I�.9���r>��^�c�T2A��g���/`��%*�Q3��۾��i��(U�I�`C�U�uϵ�m�\�^2qw���1��H�I�W�ۂeCy:`q���P��f�>x*4n�(,G���9��+��4��{��F�'��fPq$�
���!�k4�9�s��gV�|Ki2`&5Q��W�-~yY�
&�H�4n!
KP�o�?d�
.��#ۙ3�uZ��~��U�a����pq/��h��8��
'��$ ���w�#H��;{�xJ����~�g�5��"$�]L��>�f��X��-'�����G��3p�l�Xa�K ��$�R��Պ��y���B�� 3�݋鯲�y�	`-�rIa�+������u��g��Պ �1G�]���b@٪vn���.�M>�����_��g!X�$����WR7�k+o˕N@m%v�=�8j�m�[U�Bv��Q�5�p��� �����Ϧ���Li��*�!jEe�7MU 86��M��::��ؑm�Δ�4�)g1]��h���� )f:&лaĵ��)���un������;��ڻ��R��ۗ�X$ųT���X�]p�8��]:죀��R{j%�fߚE�7�j'�-��bk��!�����S> p�0�++ ~�V,H��FG�9?3�k�Ю��.���>h{�Y�/��eC�Ue^���%�	����) y� R���f�թ��2��ӋB�(���]ka�Y���[+����'���hy�%�JhU/��v��>)�S-�K�u`K@!�7�5#�UQ���=�;��Xq�\Ȼ�Q�H>�����Hw�[��m�g�d�. ?@��R��s�@(���\l�!�⨗@��a:i���3�&l��v�N����Nْ�3� ��L�=4%p���P-g[���m\-E�+D�
�0bm�vݶ�[!$[H3�K�;R�AxW�i	�L��:b�l�y�}\�%�#o)n�HS�+'>Y=�5b�߫gEk�g|?&Sqm�u�GIm�Q���@̚3;��l_�R!;�L����7�^X>����sf]F{8_a�q��N~�|Z	�{V�!�]/����VB�G�8��8�Ha1
����n_���d	���`�2�d�x5��&��.���)qUba�J�hlJ�6�����M����u����d2�A� v��KDn!1lFv��@T�������9�Vҭ2 �8����q�f�����������n��s�i榮�2h�m9�7��ϓ�ޡ���.�Ɯ��8�δI��t31[��Uv7��{ý�ɩCjp���)yҭ'��ϥd:LەbD�(��֭�u�"�
�+u��O;x����l��v��}�D)=$����꾮��5<1�i4��c6�w�3�ƴ�)�R�u�_��ԛ���,��-ŉ�.�W��kx]:%�vPw�nU�(sDN/d����U����_Å�t ���⤥�1]�i�$�� �0fɧ7���`�-L&r�!#� T��k$�\�"�ZG,��#�� 
�Z5H��6;��7�$�ޅ��i�șm���H�6�Ǔ�X���|�j{�Q"�3�.bvj@�!|N��[90Fb���thR����݊�ճ]�
���*��"���"����D�rx�K��<�v��wV�NC������D=�M�|�ŰJs�Z�Ah�D9Y��g�'�ȏ�9��//>h�	�z��ah-�^�d�࿃�����?X���M��[��3�ӛʔ=����	�<gמČ@�.3�I3����ʞ	�*α���Ϝ'b^Y�&���9;Y�COK#��f׺G�hg���{&�*߰���5�t��YC$�WԈ�a.ԧ!�^��2Q�{��/?>)(=��*g��������Ĝ	N�SO�m��R"e-� ��Gţ���It��8O0���P�C�"XV�z���ɵ��3꣔�?j۪S^g�3��ᗠ���v�)��v��+�Q6�^���b�IX���3�����p��Cp���ؖZ ��9�^���f��n�������6k�u��<j1��H��G�s8fn�X
*���"���G�o�C(GK[�:��4FS���<���r}ۋ�`�-J�Ŗ�3)WC�s�by��%z�C���gX8{
!=�X#�
3� E��_�E���cQ���#O�i��j�����q�M9�Y���+���t��E) ��ʤ�j��eRι�n�N��0�H0p�.tl�j���j��-rx%쎯n��e
��4��Q-;�c�{J��ק��Tf�>ƈm�n���ڴ�c��_����P	�`ggB��5lթ���s����"U�Zs׌K�	������i���s���pj/3��ja2����|::|͠ M	��V�q�{��b�i� %�%
�j$"W^j�ו$Q0�h��7�&@��:t���Ϧf��Qb_�:$w/�*��sǉ�,��/��h�P��'�u� 6�'d��ԙ����A��6��W:����V�����u����Y�M�i��y�"�,�=��jH0'c�}u���{�b�����NO�)��u��_�~o�OX�~�\Kc,��(���-lx~�ud4/�F�;ݮ៯� /9��Q������$��QC��4|���M�U�5�*��vHʂ�ũ*>u�{�P�0~t��o-�Dr�cw?4c�kP��a�Ee8�M)~�N�`g[ڈ��d��A���@va�/��0g� �,w��yIA�=zd
���P��6�	x���"z��R��Og���z��p��k��FB�*��v��B3$
.��	d_''n�}���"�I�}�,���Tp/���|�v�PD`I���Q�����E� S���Anj�C�/��0 w�A�s��[��ֈ0Nw��[U���Pe"� ���9DT��~�P�z9�ᛖ�`����@���Q�7�5*Ȧj�t�C��M�!ǤM�((��.$�6>B|��A.�,d���37s��3�e��t�xi/}n5��F5��қ�򺜧7>�:߶Hx,���&%��Y�~�g	��W��Y���2�H�^ioƻճol�	 +Yj����4rK�Ql�={�
�$��H%�;ח�����<;�t�d�0����&.�Lv���(kuH4���n"U2�a�yKBe��'��]T�?T{_ ,�'��p|2/�B�"�=�1�ž<���w_�5���o�G5�K�T���b�?�A���3.�!�,�^�:��L],���3* ��mb�I�����:���Sx�u����dr�'V��T��X"@cƸ�j��F�;m�|T��v�@H.�WKgF���C�lB���d�A���&�6���{fT㹈-}�oc7���Z����N9�,�쇇K������7z�w����Z/���eJ���P�7:�,'w�x?e����{��s��8q��L��*n1�d�lq�&|��H��"
Yȅ�b��k���$�c�j:�����mS�������>{ET9�1F>
�����x)K����x�C�I���	��U�4�6ugy,7c�!����Q�*�����T�����wX]�)rZ/XvNC�.����V�u�Ϳ�i����f@�7ՒU�t��-�G����vɌ���N,LU�:S��c��.R��vt�uuZhs�?�G�w]�+.���#�ǫ��ɠ��VV�	����q�����d[|�Y��#*�l�f�IlO�@��|iG���;o2�p2� [6�-*�6�ո}z;�R����u�3��㒹z��r�AoXŹ��J���.K�,�Z4���*��|8w3K���A��3d��̼C}���V���Gȉ�E�s����������~߸������;��o�^����Q3P!�E������r�+*�]z� /Ǚ��&��	.�$�Ħ��@����� �iʞ�C�A���e2S������%�$�TC7���k�f,o��l�Ͼ�D�؎fP�v{҃��L�!�m�84¦����y�R�Ǯ�ɥ�tj�a-���B���~:����ZW�|���.36��-*\���#���Əc8ؠ.$I D[��`��%CH=@O9���f��i�(b�T�.P������B��q���ͥ��V�?� o\��O)P�9E�#��7�_H6��жQ�.vH*{.F�	x�;����m)�Qe���a>g����Կ��>2�C�1ZK���Q�sJ��,@a��19�k�{�)u�\�ǝ�{��[�q�Bw$���[ބ���2Z|k�yc_^C�º簴C�4dd�{k��NNdoE���\W��my;M)�@%����&m�~����rݖ�C1_�%5�6��~�Y��g"XJ������������O�z݃�Ƞ��;o#/���h�(���2���DUVPɒ�XHI����_�;=(�O@�d�����������EB��݅��L?�gE�[j�KqҢ,�v���|�A#�*�������_�j�E11W6�7�q�a�Z�,J+��P�\�~M�S��Ѹ�s��},R�����V��DH��!�B����Rx�%.�� !?
�@��TLS�J�#�$�~��̑L�*pCB{�z���n�,�fϼ�n=��7�^�ƍ�N��A��g�����%"q ^��"}��Gn��_v�3�u�*gk��Ƴ*�.?�^��&/ ��1�A^
��fC	�.1��6µ�Q܊�[��1�hnܼM�DP��%ϥZ�Q��a@qAy�	
�q�E�Jmo"I[B��Z& �б�����Hڣ	���>@����-U��AH������f�o�Z��\��T���K����|0$]���YkƁ�H���*��ő�4fw��OR"8�C��zO�N.�̇�N�M��4���z���SP�(�6驸H��S2�˜�4�<S�j�
ؕp��
$>-��cN��T}fz�=>RS,`Qe�̛�ȕ�1���|���%}_|�U����>D���_�dKffe�,ފǑ���y₠,�H�]j�a�$t'����V���>t�u.ckF�bw.�x�Y�@�*���,-���'W�t��E�� Hy�!��fd���7�?�a.1}��Ycw��=��k��.5�1FĀx�`J�muW��J��4e�A�
��@���MP
�7ܚ�`���?�X'�{�u�|1"3WnQ��m�;Q�E�N���~���K̛}�t`�o�N�P�ԣn\��ٻsR
���tKc��f���J8!~�����pA�H8�z�+d�R\菮-�3Ū���5Ћ�J�Pc5���f�߲�{z��3�g5�\6z�!��U��`͎�lnC<��
?MӍ����cxn.8�ۆ��f:\}{#Dh�4rP<y#S�L��`�3�#T��7S2� z��9~�A�2*jgQ&�
]��Fs�͹�� S�D�E܍��a��; =�8q�AVFx��#䉕a�S`�}�j������xf�8Ԝ�nܢ��� ��̒�8㞿���p�(�=�V��Y���Ψ>����!6k�O�E5�N��>��@�<,��܂ �x�d.�8Ww��qY���V���Є��V�����==mSKx�<�6�e:�<~cU�]�o��wm��O�M�|����)�jc�e�:��M���ZN�ALw�����o(��b�+#h����5�u%;qd����>,���Ѝ��@�W9���a���d����.=F�d!1�_���,vonR/w�d�(̑�(�㓭|{��u�cM� ����6�^M��֫����y����Xh%a�����jGIY
@����>yũaBEN{� ���-�!��;���r���� �
~�y�)b>���u���`�BWb�۩����?�r#Bҩ&9%��֌�A�z���m8�3�.��L"���-�I)M�a.jl"{��"P�cM��O%���E�|Q�qď(˵K�*ˡc��؍�Χ��Z�=����b��hr�f!�Gd[@WBO���-\��!�Q$�J*k԰����UDaqFǪB�n���D�$6������Z��f:�_�IJ��,7y4�ی��D�G�:�/���a��g��G(46VK��ר�����w�>4^�ë�ź��@����!�@���)K�~�f��Km��K���L��uR�5�"��[�	{�_����ٕ�o7�z$�������?P�Mn�*�f���~:�9#"��GZt�Gط%8�	,!jN\x�֨�aĤCz�u9W� %��o)9��)\Rr^نhe�U_�\�;�[f3{��E�V���u��N���ad���<���J��kؚ��4���@x�?���t�A'S�|����	�������S{B'�"h��l_�*��a��N����;���+�j���9J��/꫿�SFTm�t@t��6�Hʥ��'M&l-�� ���XÅh��ǩ������Iп/�عs��:�4��լ��	K� :{����5��z�<)����jp�mq{���t@���>c��KK��C�×���)6M��>{K�h����K�Jd�e�vr��,c��}���#�����W�`٬=�WD\�p��KJ:6��M(�G���J��Ea_+3�����ȆV|2�ů��JV����"��-�aD'�E<�tJRY��(��	Ġ�iݞM��z4-�[�6�?r��_�D7�4Ľ�hZTKaI��Tvaü��WHm����#)�\�	]��%)̑��QFu��$�qup��M1o��ڇ��/9�H�-�\7���.�+�K��w�jw傑�3ݸ������a�Xz{Ɵ�� 듹��̫_�{����Ϝ�Tb��:5]0��'{�A����V�<sD=� l3���{zZ�Y(��>.����n�1׃�N�9~����3Rj<��.���{��G��KLG D��ѐF���D�eC�ŕ>S�	��}IqY���ӌFǑ�x4��3�0�7Lf��K*�UZ6boT|�y4�MLn!�{�iFG�I�MY	�!��s�,���,�6&n+T]��{%%Ja7#M�:��H�lԀ�"<�ߩs3�0a;���u=Uغ�����q)�k[k��1��X�%�|B��������V����F�g�B���ʴ����u�V 4������Ԅ�*wR۲F�=�궿Ac�y����,��	���Ab�7��j>�;��R�Zy��ŏF��� �h�m%Ävnc�!,�m�1)�7��x��:�Ȅ���qoY� � 
;Wؿ���Ui%9����	�G���˹��i �ُ�?S w�l��Кs[��yԐ�(f��ǂ.0��`��b�!��?@o��&�yk�Eb^��f�ld�@<�#����x��QX���	�?�_a�т�[f�(_?��|���¯a���2}\�>�*��aB���k�xr
��[L~\�|<�+#��i�fXyu�a���Џ=��c���@�U���v4��`�^HO�,��O`GS�-��.-nR�)G�X|�'��� �oT12ɳpTt���ߘ�jn2G�����X�_���ܵ�������$�Z�����3��� &�'��a��=��G�)v����m�����1^���	�*$�T��Z�xJ=��9>�����=���=������I�-���%�s�W+�祽M��O�J�<����hH�A��V���ħ8�t�"���8�+����}I_C�֚գ��R���A4��kr�0��������愝�շ�[ac
����y홿��<hob�u�wP2m��F1�yu���8	����R�<H��5��ў�7���X-o�=����9�_�H��U�-sə̞Ɋ�)�[� �Q��Ӕ��bw�`�!KN5#<�Y��S���`��)j�a��e'�H�c��!BU8�"�TG��'o�p�C�x��1���xE(0/�p=�@@Ç����������spr22d�uȎ�]c��d�}�fH����˄r`J1W͔Y�ꓮG��ͮ���ؽ�3jb%ǹ�NV>�N%�Cܡ�s�A�ּ����k��Ὕv����} � ��!���8�/g����1]�K7�,t����?�\�����7W��ֿp���� ;_y��C���s�E�h�~�s �/�N돥�{e�ߤ8X|Y�74N��e��lW�%��%I��'���c��42���W��>��b��T�T��Z�8� �u�m�?T+;�k��1�Xр�\OD�bB�r7u�p	٭^&ǻ�]�!�f���\4|�	����l�?�|;�ZTr,sv^�Wf�u�.��o�u�v����L�fa�N�t�-����Gid��ҝ�=�ٮ�ӗᔦ3	b�; �t�6f�Fǆi�C� {��¥4ݍnlQ�S�G�oL0�%yX:{����a�q6*y��/-D��3�>� �9)�!6�h㞳���⾯��o�b��01�klC��uф~���[��t�8x�n��KO��{��b��}�Zv	�	�G}p�
��5��?�=�x���g�͞���4��#��:�~$�9N~��ó�QUE�g��'�J�g��>:��҄�r�s�"g��7�x�uY���D���G���b-o�U�)	��pǈ��t��̗�l+�C �d
�%�] ́�f�tȴ�;7�ڰ� '��4��'E��H3�EE{���}`2IB��D�m����T����B�<�����,��*�3HF�əg�{ �� �)��W��T�1z@c A�N�l����D�S��-���H����S|� �>	�%˛A_����d�k��v�co��ͫ	O�Sde��0p����#�.vK���t��n�bW<*��~ӳ��r�Z��d�Ȋ/���e�u 3m��'�?K����w~��p�f
�^����6�lǼ�Q�!v9�ƾ<<�4~=���@1[^���j���r�KGy&2�U��̼$e^�$%l�%����kTO�mQZ��3�蝹��hV��W)��*1����(��%<��v��zb�	�}�")Z���0X���O�4�h�w�<��E䅁�9;&��A�̳K�(�t{剢��w�@�$��>l�]ʔm����Zq��w���(�Xi��0 W|���ޠ]tr�ɴ���m��Bc��XII�(�k�	��Ձ?����:q�JsX� .7���!�9Q����f�����R6[����M�^��A����2D��Ԛ����
�-&�V�^nn�J��	,����]�����o�:�	� 9�0Ehfw�U ��WMw�ѹ�Z+��� �ɻ���\��.��b�5��/r�.
�{�yޔG����أW٫�O�U_ce��O��/������!�T��� ���,r�T�Q��$���{�v%Ğ�1R�I�v�N3a�c?���j� �w��Y�&��o�����l`��D�ܳY9������V��7��(k��h�}W�BDB���RG�4��vp�\�B�#��MsD�@/<0J��Q&>��"{�˕b�k� �)���ky�!��!+��B�,{���ua"<�x����X�q �M��`S�8�ƛK�0��J9��7/�rf��K��c*6��U�\5��ĀYG�Y���扌p��I
M�*Xg�����3I�봿 ����#�(�_O�٧8��?���{䃞�	����ZԱ|b}wa��#�D��������C�fȂ�K%Q_�T�4gӒ�u���$�o��yF:���m.���	'��y<:�$ē�--���5	�����w�7UU�����	)Q�d���%��8�7�|����ò�y͐�O���H��xGq!�5fuЖ�?<�A�u2Bl�)1�5 zR'�P�,��)dr|�����"��Ŀp�ޟ�dSN1���bK��8�3����I�tkJ��a�O�F��r�OD9��Y˭?sUT��޴���叉U��X����Cy/qWK�l��b�aq��4�	�$�;n0�x��!;4:T�� `�fe�U�mj��,���krr���︵p�ǊF/�C�N��OQHy�wC�\�-U7�"�ȧL�:z�D<��Pj��@ *V�Ho#B<מ#r)�~{`���@xkŋ��h���DX�PK�Fٚԅ�-Y*a��%� ��3��R&U�-9�N���"3�>>�H<T;Q�6 ���(�/@Q�a,qz�&���^נF���rÜjvҨk|n�,^�l�=E��nx�U#:��:�Q�k�y�Ƴ�N^���}��9}*Z�
�i��}L8�<�T�J
9��i��Q��
%�-֖�b�Y<2�)�$�X��r����~C�����q%��6�'�v�G�ZG�	���X&�gS3d�9��|���'f���D�W��<��TLSD�=�I�����Y�=%���J���ӏµ���	�ؘ�5�42�1AS��i���m���O��ٶ�6��Am�W�o�~13&�z)+����`G��?�� �Vv��6<�x.~��9t���l�ڛ�̗w��Z�i�x�3^��(s���o��k�E�fR#9���J\UZ�[�� 5��z�&Y4�A�T�A�3M�7h/F�b-��<\�|�@��%�'zD�"͍��׊|��+k)E�WUW�/���a��-6g����Y��j��ȢН?��*j@����Oin+��bt���4����
�!>�z`��{ýsVO���Y��A�����ʒ�C�+��,f�r��v<Ǣ_�_p-؂ #��+E��\Bf^J<����/��)�.u�\ѣ���R���Q��.����&V�<��֫��2� ;[���EU�=�l$x���S��0@x=�h�i���,�De��צ�g���}�DDE&�c��s�������/k
��E���]������=�f>�DP7�f��N�W��ї�p@�u��HuJ.�߉��nl��SV� �FQ���5!4�����-�Bh�{>�O(����dAB-����n�7֝Fy
� �V�5ö}7�:jF8�<�O+�0�|mo�v*�,���8������:P���4�;����Rq�8�*�!6I��<{�J�k��^}��$��+��_I3��(v��hG7���;���T��P������	��3���6�-��Jvd~���3S�����3�Sd����׬�P����y���/�+Y�G<���@�F�t�_�%�K�|{R�L9�k�:|w4!�M�5��r��wc�k��=�>�}�E���ͳppWI�ǎ�Qd�w#��A�{��R�7V���-����,�y�|sۻ��? �R�]7�;DG�H�Me,�J7��������:>!�e�ǿALww(���L��⃕�`��)3�c&��#*J��j-��L)r��[����n"ÛY�C@�J�Y&�ǵ�q,�6O�A+�R�CoLK"�	~7 I�y�)����aae�����#�|�S��h���ȶӑ���D��w���7���`S�������_��\�|[+��7�}ڦa`�`>��M���D1'_ �["s�}R�a�r��C�r� s�Щ��������޴ӗ���Qcpz�n�j�N�7���i��s5�}wx�d>�H��r r�\���'2�S��(tp��8�g 3��S#9\m� �q�΂��N�(��\v6�bB>B6�f8A�[���j6�i ?uîޙ�/��ԉs�S�n��Q���0��k[9�n�؏` �G�����~�����8N5~��
��z*�=�n԰�$y��Z6fQ���)V?�Ѳ�2�f���t�ѫy]�"�	�nD���SJ� B�[���AZ�<�����kP��e�"�1\��C�3a�xb��R��S��L�8��oX����9�Lήwy}ؖ���m���X��?��8���bJ	w����~�$���(�S�$����I�g�:�-%�IB������j�)=\lɄ�l�P����D�}��O+��H|��g��s�,^��Q�a&P\�ޘi�� c2�u�[��kr��vӯD*�;�Z@�ը��9qF�6��*�}6}��V�N�Ҩ�v��i)�"��t.��xK;�[u�یX�ͥ��$=��%h�(��#A�8D�A<�C<���;����KEjǚ|�+qj�
,�8�g�m��Y;��[��Q��P��9#����'%t[�2��%;-X�<�$�[sj�*D<.(%�tJ}�#珩����,���e��	�R�W�2��)O��V�0��mY4�s��+<�_~���*�:�����k�!���7���Xk>��.�l	Wp{��{�f����~�e��=�v	OQe�@q��w���ĥ4Y^�P0Y�GLŃ�GX�f\#��soI�\Q)�n",����.X�F��F?�'	��n�ā�5%�d���H2?��Bo��G��Y��M��$5n����}��lZ]3|�vч��X�ʕ�z����C���s��^��/w��"��-��`��7��"�Fwn����Z�&�uޙ@<b6������M75�����X+���5:]ci0H�,�{��N̖��\�1�V��Eč�ӧ���iǸݗ5f�������
��s"2k��d��Uf4�{������m�嗾,x\�#6Vt3c��� ƭ�'�HƘ D}=��S���қ7 ��ĖX�s5J�j����4IG��Ż��9�|tS�@nY�Y�,[��g���3��U'��"�O���!��`����=o����8�)�u�3�ǥ'9c뭮G�����h:���:�޺��4�o�!�j��;:5��S49P�0��z��r�oF y��W�2~����4\�\x(<�[�50%�9#m�'A��cc���~C�]gUn�� ��;q{eVU�d[�N�I2^�~��[K�z��3i9/��#���6���M��J�m�8������ؼ�9z�T��-H)���� .Ƈ	#���y!��z$=�����r��*�K�P_�������]�ȍ�{`�q�
�s�i���8�0�y�X�@v�����C�ԟL{�-��Y�k5`�n�7����}ɺ��}+i�rȥU�]S�J$���Fd��?W4?��b�q#F9��$aI�v`v�c�n�Q�
�Y�Z7��sz\�1���T��,�)��N�/vE>��+�Eр�	��"]B��c�� �Lt���L-��1^�m���F����iʽ�[��?�ˏ�|�,Z�7�7}��B���� LFf�<�/����(w�Ԉr�:Zл�1Ĩ��̝!p�;��zHm@0֓h`jZ}^D\���n]n�Q\P����v�s,��xsI$�@�bxr�"[~E���_�Mu�C������Yy'Y>�D<��3&����=h�������ݠ�鳷�����̀�b��{����l�.8:���f��W[�Rk�d}���(vk����mp�� ��!�l첽=��	o�qI8v��`�š�(SB�ޡb�RE�O��Í�@l�=O08�0�b�[�À�G�+��O:��)j����7�vp�;�^�n����L`Pu����¸��1�QJ�*�j:�A(ѫ��g�H�+u(������]�6��_d���xL���7�H�uc���Vɣ<\���Ɇ�~T�Tt���!yd�2�g	�D�c�&/�c��b�%a&��}p�Lg�� ��Ck��F���h|<�|J�WK8��A ���}S�H\'�,eH�&�԰->Bۤ4��8��S����J��]Y.���(�ʢv�O
Hf9洐׊7C˿Sf���h�4�-ڠA����AKxZ�>V
���9�;Q3e E��\�/H�;�2�$�ބ����+����5��N.R<#DfHl��}��������-� l�M9�t�	YNSA�s�D�����u<�r�����M�nrfG��4ԯ�<.��}~�d�*�v(�^2��P/���v �M[�D>�����E���.8*LAn��ER��>��촛Oi6wڒ^	�sր.u��U�y��X��/A'�������
���w)���^�c%J!e"S���ข-�9"����"�{nd��qL������� �%��&L�F*:��q�T�;�<(��yV,P���ùڑ=�*�z����#*H;�"h!6��V	��o꧁f���Q�S�98~�Nl</�y{��ۻQ�H[�cʓF�!@�%�~:ހ�*\�G@lr��W��"M4୦���J�,UyCڅ�2���X[�f��l�f��h{�2z+L9��~�ܚ0�U�wi1��8;�0牖p�P"L��~b��
ĝ#�`����ôQ���7�K{�W�^�-����?��UшU*o��7��ec纁bY�ҩ��x�(R��T*���D�Ɍy�)9�3r�I��.-D��d�kA��U^��,/)ĉŏBe���Q�q���4@<�hLk�3
[�&��[�	�����#
G�m����4|)��~�'��m�� U��f��/"�p���3!Of�-��ܭ�E��.J���<�A3�s�S1������񕵸�.���g{�lRNLM�mn&��F�Pb_hm1^î�Fu�v��.{�)��EBt��2��-[xm�6�mG����dvs�&j�Ծr =�䌉Q��{��.��sq���U�Y��}dd5�t�6��b�w"u��u��'�;��)�Ղ��z�<�������eD|�nt&��".~X�|����Fb?}H��"�p��'Ø_j?(�t�D�4�ͮ��݆���p0U���C��l�\YэW��Da�#�%���C��T�K?;әc�e�ST�T��9��HA�Ao����Ř� ��)Ia�~}��w�~@��}�Ӌ�y��X9������2dCͦcߋȶ�IW��ĩ�w�,��;�4Oϻ5Ϸ����(T�;>���|��Z���s���^ S��1��r(�hUs^�5^gn�.��%0����$l`s��\�|ZQ�my�pJ��~�/�+�uU�W1P��"��f/�Ŵ�,�-��Ja�f�����!�g��Ap+����ْ�:�`�[���+��3��T�z��$�8�՘�O~X0�p��U�O0����@��F���3�k�KR�j�<bl?|���=O�A"G8a���Ze���D�,��&�K�.i��@T|˪�ثC2�.1x�o�þR�˽	�a�2 �7�D@o���Z��t��fMvb��/��Q����\�]�{ɨ=���'�+���ݩN'�� P�9d�J�U;�0�|�v�o�=�ZX ���[Z<�A@��;���e�|��II)QKΈ��AE�6G�"��j����*��27�DG%�����M��F�>�I��1p�	��P(ߔg[�e	��I�_`��Sd�A�<�O�Z�6�S��H��E\)�s�?6�q��-�z9�ƶ�� t����MyU,�&1W�JGRi�Q%?N!�����B�'��`������걒�l`�s5c��g�Y#��V���Z�����|��'�~p�:�ż�2�U�՛�6���A�{I���A�ܾ���X�Dװ�����~�967���4e�����P��Y��W�ʍ�ckF�֐|ʙx2�<N�b�(�āJ �^�孴R#�?08N���LD�8��5X����a��/�j  ؜5�%��{ Axr��YЪD��;���&=X�ds��y�5���L��{"�۵�ɖ��&�l�~��<�ښ�iT�M�g�N��GCr�5.��>�%��^t�� � k�-.I����oR���"1Ģ)��ز3��8g�OSc�	��2��*af�w���{�&�� �]<���ۺ��#�����*��E� (��o_!���--nf�?��/�ј`,�|:ވ�M4�����7��HƆ%Z :�w�|�-u��D�'uV���T��1�g���D�4���#)8-꜃�N��Z�#�l"PV�zP��2�\n�-�P9�>�<�BFV���/�.3���g�~\�kO�v4�/��5?���I��5xN�L.h�C������+�G�'���4\/�a��QHى��YFT�jP-(|�s�6}žݯRD�7�2����c����f�P��j��`q̚Z�~���>���f3�|c/p��®I3�w	T��G�{��ǈ/�`����_��yJ�X�N$8:��i���$r1��C�nP�����g����G���a4�&>�`O���0�S�,W��� �O����ا��Rl������)��@�xN�"��w`ZO��0�kѫ����4_������t(0֩�h�+C�έ��?�O�h
��X�}�z�O׏w�9�w���R�,���G��D�#q�BT�34G��x���#]��U!%*�)|��1C���ݷ�����4c�v��Z�ђ+���u��CN>)ڮ{�y?c�9;��
�����lF�wOD8������uz� .��O9�{]�h�}�@��΍!���>YG:������/l��27ԻO(xX*�U/�jl>���6O������7����$Y+(��g����/)n��
���}Zݜ��E]��O������r�	)r���,G�G�!&0#J��Sy꣎fx����v���M~��YB��;�Tq��(Q��C�b$��Jnް��!�+��V��8�FP�=���G�IQ�Oڸ�ՙ�CU{��7�0�u�	���:tR[rK�3M��X!��sbW+,�Nǀ}��V�h�,?��2G�4fA "Z�H�+��, O�L=S�ﴋ$9q��i�N�+�X���{MI�t�m<gq:���Ym�����D�/,�Q++c��H/Q��|�FY7k�T�=�0]l��p7E�7��mq��~t6}�bAz��+��CqB�g߮..�2��2<ا�<lLN��V傊LY?�mءu�EC%Q�7���me��ݸ�*�B-���Ũ�`cA)=�ɱ�Mr�*�u�sf=�l͆�vc��K$�I�t��&�M�dU�Pn,P�#P.O�k=�P�+5$��a�W������a3a.��>���ܒho��x�"T�KEE�>*�ϗ�rh2�Q��ˉ%F!�vWz��´��#*lbzO��7D������tT�H��F��]]}[ټO�ꁈ�B��]�����:��b(���{�� i7�"Z�r���	��\�s�%�r��V�5�ki;U�l� VE�dc��޿@{_E-��نv�>J(Od6s�P&z�i}���]���E�ӳ���?Gيb�mj�c�8EJ�6н�}C��_�C���l��;�a=��׃�/~�/�������:t�M`�p[b��=�'[��sC��k�l��S��C���	��Y0 �B}!_�a�D�v)�ϛkrt��iT�H4���'$��4���gڷ,��_G�j^�_��Q���z��{@��S�7Xؒ�t�٦7<֮��D�=8���X��VE�hjDuR��$|��T� ����|����e�w����Ȼ"/��1t#�`����4V��A����u����ֈ�5���
�$�nCAXϵn�ڪx�P��I��-"Ĝ��C��=�\`�"b�P�?����U�֎����9��5�d[!���0V�LID�bj��/DX� +��'��ݝ����B�7r?�Ỉ^�����UY�֑�/����� ���٦7�n+�P�c-vI=�c剖0L[���ۭ~#JJf�'�ӌ�NY<����w� @s��rZ�W��}*���xI�Ǣ��	��������rO�<�.�.��ϣn����'(�5.@H���nC�
��X��D���U��/4˚Q*NWp^^��]L�V
�2/�mQ��u�8;�KN��#�VZ4��$*NOs�6 �$�6��N��������71�N��JN�ݑ"��-�FT]��5A�2,��287O5׬�FpGX�]�$:���eG��vzFZ� ��0s0�Ź�U[!?�n�r�H���,��8U7�ƑeG�2���	�c��:z��{��<��	?He��ډ�e���Nއe�f}��d5a8�Z��3u5I�A1['��Ir=p����lϺeX|��Z��7 �*
S��I�I��k�V)�*V��KM�?�+�)�6�!�u�M��;��.t�.�;�I���ĩ���eug�a?�!��W+?�'|�`1�Rɹ;����P7Ȓ��)J��^$X�i$.�,/�~:1^� 7,) �Z�ֹ�3��#�2���u���=b���'J?U%s�qD<� L[I�^�lx��9%�|O� �U�'$W��13*���J�<��F�p�h���4�s)[�hQqS�z��ˢ9�ۆ.����C`ov�^�I���5KS��8���i����F\�in��]3}��D��u΅X���E�qlNB����_!M�/b��'��b�gꗣs�g��AMR�=�HݟO�'�A�L���G��cxVIka_0_������0��=�iGS��t͚����B��C�ũ���P�
�`G���l�*/m��q�_��`~�L��=����go�!�:�څ�>&�D1�$Z8�At�����	x������T�����EJw~�Q,e4�=�&�&���x^����gS_p�ܩ9�e��A6�^c�Ji�؀�v�O�ΰ��j�5-n�*H+���ͷ�A�p���u#�3�.x� 4�}�E������?��h�F�@��`�#�݁�7�s���/ʂA�a?U�R��+֬W����&C fB6^ɯ�l'���M:��ˌ�Y��Е��z���><��?�2��*f���z���-���\��!X\ܠV�{�����I�Z�(,������O�_xa��ޫD�x�z�℣��<�O�Euս����C��,�'��ݻ����i���N͠�YB��$�xCR�i{QTJL����������X��,I��aG}i)���|"Xīp�gI-�q?�&z�����a�JVr�Y������(EX�.q�lQ&�?�Fo�#�ih_JEVr4I��q��YK�Dg��b/E�����ٹ�N�������m@��&��6Ԍ���0�6�i{8β6��?��D���׽W�2X�0��i�8����6� J�P�h��*�;�~2#�8��e�ǅ䮖��]�s��L�!�L��ta�^^0��a@�(�9����,�B3�H.�z[v�v��ns0$�L��f�!ϼ�G�n�:�:�8�uYT��B$1��H,��|z������7���&�L"����H4{����h���vŗ�5���,#Vn���2��q��������Eu�P��ԇ��2�f�f:k�.ÊE�a�kpf�z���il��4�-.�	3D���qM-��L��S��c�����)���{f9Ҍ�1�D�B���TuaY{�m�&ۡUg$��s-�@ւȞ)쪘Hx����9�(��M��h�2"�ͪi�<���uc��c��^yY�gA�+z�a�`��7�^�d˂E��ۖH���mCЈ:���*VCmGAA5Iԙ��y�mi�,�����ω���\��n0�v�P�Ǚ�Z� S����,�a�z�'�Ay�}]��z9�����Ӳ������j�AP�'Q�����w�@U��q^ZP�r�Q0FHlOJ���.�GAZ@�C��@�� �����z9�2�>/�*O@$�c3�1��1$<��7S)�~�sgT\E׸�®�.
�37�~l�����a�j ��}ݑ+�4��+������֣]����P2^U3�+�UU�P8p���V��x�N&~�m6q�SKG��.Ҥ[��m�1�nU��P�7���NPĸ"��cRy2�q���YL\����F����Q����`�&*�I�fz�8IE���%��_�,��%�v����؋�t$	�^rܖ%�`�?O����3��tLy��k:&>�8\K�s��GD2���[�j�u����i�����X)a�{R�}^�M�wU�S�3-���A_fa�!?��p��+�h�'�4��`P�9�zg�i���WPZM�r~�V~�U���/ w�x9�T�/^��c[z������We)u���ކ�~$��a�Y��f͓
i�f�z�ї=��E��5IƦ�F�Q2	�<����<��oX9J��5 *',Χ�zM����+�U1�	OCi�����]�j�Ge$qN�������Y��Y>ȓ����,<�(�*�S|��n>c��\�2��2��y�"1&5A�#R�/f�V8H��?( �ᘆ8O��Lw+~@r%�&����c��8�K����*���U���;���2)n�����{s��M���M$�{�b�)	Qk��<��"Q�����#�^�Ejs��oc`O�$ ٩���9]z%W���=`�[Q�ȋ�\�$޾xw]�R�Li�� c��Zw�$'{��Ȼ5���m�fc��K���Q�]9��X���Q_,��74Hx�"3��������t@hl4���Ғ�`�SSeG;�D�Z��{���.��'�0 ���u����~�R���������q���"	B�X^���`D�)II̟2�R�������߯�����d���H���^c��aC������[
��fn�r��|"E����f5լ(�#�P:�l�.S�_T�)�E-#G�Fl�v��"�E�����HS���^5��{V�!�HT�^���z2�/Q�����1�"/���HK0&��A���Ԭ@�
���{)�M��
������%��Vg�o�1�_/?��Ib(�>�����ԅ�P4����וX��	����Y�QM���,bt`�X��_�s$1#��.vI����"`�zO{�u��n�io|����ހ���I���q϶u�^=�յ�#�T��H}��]|bea��!J�i[J�QY�Ļ�h��,#�	M���Ԁ�Ȟ��.BԹ��~�
�S�<Ʉ�%I�R���H\�������-	�a�|V�4B4j�g�2�g���#T�ֳ^G�_�1�	���J���g�}`v|uI�)�
5z��8�ɘ*��J������_����l��4ܨE�oA,�N#T,�5t��flOᗡ�6P9�)	��3����7�"i���������4�q��,�N���\�~L��x5��=�ZA��su���T%�_P�)zֈ˔��,�@B� o��k>%oً�_�)�m��{�V��4�o*�6���u#�����?F�������@���]�5ª��.1�%������A|�L^��� ��$�����ЗW=e|0%^����́E$�o�-����ٍo�
�0ؙ�Cr"mT3���q<I@��us�����kU�Σ��aux'�������U�Eѩ:���7����)'������8֊�r�O����=̀�7n3kf"<�W�;c��Y�N�=V���]pf�:Z�e<B��:�����HVn�2s�
h1�;�7�;�t�k�NR�Sot*j�r_�a^Ǐw�r����-��>l������N�x�P��[<��x��6�_��D��siO;q��E�BA����H����y�M9���~0��fK�Bd�Ts������	�q�l����=z�1X?"5���k��SZ'���8��ֱV�l�@�S�U�|	#����M�R���L���֬{_s��Sv���E=K���]�AS1Z��� A�vj� _˶k�Т��5�#�.��E��Wܒ[l@��P�2�Vij�݌���6�~뭲��E)=7�6�[�~�A��V�u)#AyznJ��}�"�o���$T��\xb�[��{=
m�8y�#������>���@�VI�r87�
"���l)��Lض"��>�∵Y���.6��HM�Q���M���݄�^�	�Q��'���:<L|��?����� yk���y��US��@����|؍D�N���)�|��qz�Q(2Asoo<�aN>esmܝD9�^�%�4N� #��i��
�q�]s'�4��0�5��D=г��]t��ǄK��_SA�����E3NT_��o��-�p�wT]�n�L�kr��ۖZ�3/�c�������|����4�2�O�㶃�hzo$��m{�eOo?�w���[K6S*�-���/.6�*��܌����逳�̻�\G���0�@����Ot?���b0�L ��c:��QЬRX
��vV n��#�>E��D.�!dP�\�"��Ϙa���B�H6 ���oG��.B����s�U��y�T ��������]��Щ���<̼/�_��i[��c��x�d���h�~�_l��pq��V%-�}DjL�Ţ5S�t?8p6��鰷�� ��>��A]N��%��V��!�e~̟I��>�F�i�1�ҲP��]�gqi�jrr$�ze�"p�!�/?2���p>�8�� �8e��4űqSm}jB�]�})}>��[-�oPy*��Ҽ,���B���HA���[�+x��,&��n�od�) xo�����ޒ�\,�ӭuN������CP��#��*�CZj82^�2����E|k=}&&�=H#ۃ�D):tI)�1Tk�+4Y�͛b�x�_N}r1���E\��i6i3R�(�m3c��Ϩy-�1���痓�����J���5�.��7�:�g�YR�T��c�K��u]*����ާ�t�qE0��4S��-p���'����~"XO�������*�P{�m���u��_H���18����Xe��^�U���'ܠ�7���]_�(j���]M�9�S|̪R�6$3�h+��Q���=2����U
����B���ז���<J{1��{��ݹE:�[(bc��������P���8����ʂ�����H����3W�2h���.Z\`����,d�FcQm<uC��K�	�_5�뚍 [�mȣ՗�cЛ�2�Ϥ�:&��夬o��&4��%V�
s
��s�7QNǿ��� ��Z���o����tI�[���^�o��S�����XZ�3l_QK�����b��7s\����'���+���r3-f[���E	�Qaq�T�F��7`��|�5 Wj0>�UB���.{Q�|���s䕳������v_�;|��#��������x��K�G���O_�L��ú&�"�F�R�?]l!�%��߾#2 ��Fٙ������� �?����+��XDyFG��ws\��W�D���Y����%TM�_ ����A����݊:�L�rn��F�Ӭ�x#�%�p���&BUa2˦g�t1�����D�%SKᢷ��.���F�l�OZ�wt���\BI+�7�J��ƪ�Rz�R=r�bE��� ħO4������I����B�$�6��E#��k�A��|ӎK=&Z�f�A���)^1�6�ˌK>�~�,#o6<p.�A�ٳ�瀱�b�1��ed�8耦]����	e�Q� ����z�}(5T�l�f������.���s٣ B�^����a�F�s���՚���'<ŶO��s���P�xj�+��� Ҕs���0�Z�鍪�;.�L�;�~x8�6J�ۨ6[��V���gg�6�.u�[���j9XE��Wz$l��ddE>�n	� r*��;�./2`��&�B�YG�%���'븰D`9s�F�4`9K;z��2�S�I�EF�9���ʃa�$����3�X-3B(&����*���M��l8�;;�Z���#��R�O
f/ێ[�P�Fx|���W�Z��-u� ��)��]�Z�	o�b��� �>�*�<#ر<+��
Y<:�+0]�-�B=Ն��d��+]�󰖙]N��C����`µ���}%=���v���N�IU-�����vJq<L�p@&(��Z�%��z0#}i��`�0Q-I9�^_[��ݝ���OZ�¥[ J˒�����4l���v5"aEc:���hw:&�$�o �5�7���(�>q{;�+N���nz���H���F�6K�,� `����� �@�w =O_Ѷ^��8p��t#啠�Q�����T�NΧ�l�����LYO`���Jj���� 1�����T����}+&u�,0ۦAƆ�� ���3���0#��,���˕��g��L5J��=��a������T��8�i��2�I^=}�V��w.���o]�{|�8�;<���������yp���������)I������H�_ԟ9`�ߎ7�<n�-��ok�_
W�SiS�^)� Z�)�Rp������;��1RO����{,�+�]��*���5
��%
�囮u�Jv����V�,	�.
x*�K��m����i��}Вzɽ`L����5	KB@ƣ��6����A1T�,��}�#,5aQF�w��o)u�]ߤ�������`�,�,��t��ҕBMY��7"0�y��+2�ۦ��U�����,�;������_���������4�����K��j�a%f�;�yrT�i�)��ƛ4���n�<Dq]�Mk�gc�-Q��^g����_��Elqh6�q�OF�_��8�_�ff9�eQ	/�泇G���K�X(#�m�P6�G�m�笿
�O��[<R�>�ӟ�D�{�0�q�i�T��.�>p��"1)����6����k"�)�z[���6��Ѕ�2T-
��@�9zVl��Z���f�w���JeTs���c���nǑ�_?I�kqǚ�T�])�	�|�"o�&C8�PH�v���xK����+j�L��!�ō�5�����w��؜IE� ��2]��e�����)�	~�h��4;��'�e�Xk�E������:9d��}'�R� ��Q��Q��?���:�E	�8���n�$Z����18�9�E�˩��zA�N:�.���1�y�yuZ��!IW��c�떜��w^2��N�uo�4,8bt��_E�D�<��^S�A4RnSc�u O'��T`���ԇ3߻,���$���h����끐IDL�=v�s���X��ų�?��r�(����MrEVf�Õ��t[U�b�d��=ivE6�Z�
0c�|H$R_&K�V��0� .)�?mDny
����~��4��7ʂ�'���)����y�4�d�k���L��@!&��w
:���5���w����Bn/��wZǽ������P���̢�� /yo�{�^�2)2�m��wN��s�����7q��:��о��&>8��M������X.e�_����c,�Uw/�|8�)���>:w�xiTS�Hikn=��pB����̅7��`�^q,W����rk](v1Y���_�����_o� a�R�7a,[ϐg�~�&L��x?�S�(�FDJ�Rq���"S��V��agU�.�'7�ߣQB�xk�'�AN[�P&��
����k�2W���{6���.�RZ�&���\�y-��6���w�7��-JQ�V����)�x}#"�N�#wf�al�J��tߌpd��F��%Grw]H�m�D���T:9�/Jy�\����D�kpT�2�4~-�% J�r'	�z^�i(;&8�������-�&$-ҟA�tS���Z.���R�vJSS�C+�d�og%;��^�A��s!��U�߆FX���1���6���ӝ�^_Z����pk�%�!������Į$�;f����ױ��t�k"�3%8]��1��z}�l0uw�wtK���0NO����P���B�J~�mKπp&	�Z�[߲�	�װ+2�gE+��ʽeZ�	u�3-���c~��'S7��<�t�[�A��1׶=��m�[|�<��Md����6�	�)ǲ�,l�ك����.��wg��a� �{ 9^�˪)gS��|���o8|e5�^�d�!uJ�W�Q�I��g�m���O�#��xFR�%��;;kt�i�\�_�BA��IM�T�!���NRWy�?��X�E��<�9
�J��4�w &U[�¶:�Id�L�A]AF��m�=\��[�Ҕ��s�b�F:���k1 }+���\c|=�g'f���fB��8��Q�)��W�!�d$*����5}y��3��I���S����"#�X71t���D�C{�-;T!��`6�e,x��p��I�<���)�-|;d�z�L(f���?T���f[�i"t�b�&k��9���;�B+��JKU��=I��h8��[��߭�,)�]8R'�7���Y�%�I��wi�$���u����#��1�S�Tݜz����TG��q���M1}�<K���r�$pE�[�����U2�9���n�9_lG]Wʲ�X�i�C�;���ߥ64�fC�ײ�֔�ws���5��Ǽ%{[�������L�SUV���w����u�TJ��g��ߜ����5lծ�t3�"{i�s$�$K#�4�ך+kǚ|UF�$��a��:�h�:�[����I�yD�J�VA;#��[U~�v��U�2�&��%Q.��7﷛N�t���;��D�X��7wب�Q��U��!S�����_��3�;�X&��"��haj���k9�|���*mQ�����������tPOA����w.gG�=�j��M����<�u���U	�}��AB�vP�`T�������T�b:2N���}��i���c"+*������=��Е����騱��B���~E��%B�yG�1����`-��x*�j��·��_a(�U�S`2f��NC1�_b�Icb�oa��������!0vs� ,���*���Kۖ��S�3��w"_���Οn�K��;���j*�7�Y��� ���Ć�P��0U�=Km����Ģ٥n�H��\(t��ME�6���rsP��7�h��Ev�Զ����t&Y��}=�|��V�z�9�6��z��<T�Ȅ����=���#�T�>����B���#,�gw���^�@$��%d�.��	0��"Gg��y��4�%�Vfc@�8�Hyz3��q��Zw�� z�:tog|�����N#$w���]��T�����ʂU��!wWu�|���{Ʃ��J���je���*53���̚z��>S�з���i�o5�0<� �������{zcc�%�ۼH��B$���B�]�b�.���sv׊��F?�?���������ͳ�T;ޡ�����/x |C�qgu؉̻����R��:���Z�|�涣�~v������?p���+54
�{�I"�ik񠁗$t;��vG�Y�ּ�Z5���hO�S�o��'4�9�v���A�����k�c �0J���(���1Iwfo�ψ�ؼ�][��Z����#��Q�t�S��v�Qx\=���#�l{$;ˢ�ޒ_Q�\-�[�z�~%=�a�֭��U(e�*��D�RP�Rh��'�t�=�l��S��6�H�0o��G]X���ȈLT��r��?ϴ�j OE�k��%�%����Y�l�G��)��J@'{�?�Epo�|���GãD�^����8ѡ�3:\�
���`W�,ܓb��(s~b��h_�>p���>t���*E��J4�*7�ζ���)��ml���n�2`lW�|:��̀��ɧ��,��>G����5'�Y���1-tϩ�Q�gS��@W���`c�P6}�d͐�՗�_�B8'�y���ub�:iT����d�Ϫ��h�A��}��f�0a���Z��3wq�G�I(f��~_r�P��7j�1Z(�$��y��ǯ&z{Mnރ��.R}���w>��/ĵM��8n��&M*�֣�=,�2�@OZ^7���`^d�½� ƫP�!o��FY=��?�"��E��IUj�9������:T�k�')��M�!Q֙2ʹ�N���є����o�a�9�'�H��"����L߁;���`��2"�s'3h��J��~0��I���e��y(��5�� �c'ɮ����>)�'\���C�IE��8&\S��Z6��z��C盩@WU� �D�}[�>���/r��B��kW��7���7k;}ܡ2�}��0Yn�3&Q[SuCB)�Qb�8
��ٮ/J�#��8�Oc���?U%Kf��>������k!Ny/yS�����<j��Z2��h,t����Z!/핇�Q��9��Q �u'f��_̢���`��yC�x�F�n_&���I~3Pf��Q��k��@`$W����ݔR��'���Ez􎩗�2
�� ��m�#XXkH�lj�'�{�`΅��4�!�6�� ����Cgر�[hg�����Vw���z�:��1'��:�bhgnH�ثý�m�L�@V�8�b�z P���Tdw���L��!�4���*������iH�+��EV�o�gGq<>4�R7t�$�z�<)��N��� �/9&!Z߳�ƥ�V�i��14�n�H�d�¸2&�_�X1)^g2}��
��5$��8�d]�w��l��\�%*�RLH���۩b6�~����R<I����, ���蝎��+HT{�Ӕ���u,�:�3���8C���Ԉ̇,���vy�Ϗ	$5E����C�
�>� |?�Wc݅a �dZXY�v������d;�i#�I��-��m!� �%mȰ'!j�3��}��.	��,jﻁ�@X�>�
��f�0��4��uN�`@KX�uc�I���i�fӒ��$(�w�$)8M�RxV�g͙�24�F�&���M\�gdd"�z��Yf�%]�y<�2���㼥�y�Q$n\�ه\d��Q*i8�����q�N�eY�E���<�Z��Z,+�[e���sؒ �b'~��`�U��2��!�>+H�bТ-��~q>k�uPK��$��D��͏�0:*�$�|�4Z����B�\���+�`�qSZm3U��Z�31�!X)
ҧ��,B@À۸��h�����B��Z��~�$k�, y�)Y
�/�����ؤ��b�ׇ�<��*\N���P�~�hu��?_&D�"��s$�B�YH�O+Wx+ ��2��Q�5��ю�G:G��m~��Y�,�4�hB �	>a�k�х�VۿN�-,x�Zma�5�2�u/T_���(��J`5�Ј(��W���hP�xo%��(9�|~���z&n������O��(C��=�ѩ\�0O��M��g$l�l-K�*�Ty�h��l+��xDS���n;�w-[���i�'��bj�l0����i���3��~72+��c���Th��W0 �Jb�=���NP�
Q�Dn���4��t���[�t��7X0�M�9a�/Y��Eם5�U�,���4���u�6M���ȅ�φ�)s[Pnr�kN:}��F�a���Q��rE�)��
Q����B����Yc"+�8-�����VdA9����Tj(v��^�� |��U	48�<����Ѧ0*%���4%$D�7Po��"��l��zE����d;nWN{��ԏ��u�'�\�L�1�;Wh-�~�@���� Qi��Z�yP}n���sE\���i�/ܢ��ZXa�W� �m�M���p����R�~Π��e�q0#[K�#g�؁��j@�i�2R��I5F*
���'N����,W�3��	���*���_S���e�e�N[�D��Ƶߢ���<N�	 (R�vC��N�؈P���*�zgQ!���ߘ&i��q�v�QR6E��_4����]Gg���%ʄ��F2]G�C�UV�=���.й�"�R_�G�r�D�D:,��Q�Eb����S�nK|�����b���H8�A.��ɸG��ٞ��R�S��Q�)���[�����e#���@T�D3�Sۂ�s\4x1��G�X���r��isV�fN����]�(�O���l�Ua�O�����B�����o~��1�%fL����k#x����B���*��<��z>a��BJ,���?n{p}���Ez<��ؤ��m��wL���)���U��;4f��/�?��X�ܲg�<i��W�j1��'�_:���L��� ���.��B�
A�`�=���3� �!��L�1Z6�ŋ�p�F�ʅ�pad�B�j���z�W�>z5_<��1�Y�|wA�Pa�`�2P��6
�����/o���f�t�z��.�oY$��G�hSm2%�^���ec�}KF �uy\?��>���r#���!�v��C��
?!�t��Z?x�@��V-�� AK&��^�O�{��9�χ^�ሉH|���������p�:������4�X��G@	ғ��0���pm�L���P��^���F�$��-��'/��S.B�<��j^��7�Y8
n�Rt(ڞ�>�c�2ޯ�w"�G+��'�`a�F��t�� ܟ����o:�G���yO,�hrCh���WM �j`h�hw�5t.�X��P��U�妏A�|cM1����]�X�|�����W��;zPGs	����� Y�7p��Nvw�XjG��J;tjkA�I֩<��,G_��-�p7��U�s��®Cc)�X�Eђ�%oF#^3Z�՟�U�L�@{$%������1t^������̛oZ�bNǔWY�Hg>l�B�{�@�S�f�^@3ˌ4���|-��lKr�%MX��F�a|T�uBp$uS��"~`i�F�8�Z���H�N�I�*	[�f�?�8Ta����P�g�����H� �?��+�3���
�9LHH�i�8��1�w�g��v�^���zMz�ZNC��艹F.[�t27;U3~����p����͋w�4��vy]_ur����;�B���VF�(�!c���u�c	.��/!���q�o�d�^�M�WZ�W�fڤ�vI�����y�Z�3�ڵ��5[;��Sc��N'TG:>��?�
�;2��q�ΔG �
� �����	�n̝�S^���_o^�`@CH����	��G)�1mo����|ҁYJ��MïR�*����(�+��� z�D� g<n�o���n�3? Z$e�uJX���_�k����&�Fy̝�9�`X���*�7�(r�:Yx�ݲ��5�z��靨����J�a~���C�]�U§Ư	�7��G>:t~��!�	d�xI����	^���j��T���uT'ȩ��Q"૭>���d�b7 �w5���'�^�x=~��3�/�>����Q�׆x�K�9����'*d����c���5���-GBs�]�:�{�u�� H
mfx�f`'����aA�,��*��p�1B�L��J�Zzɳ�px0˷�G`��>Ш���ӏ�h�b^��48p��i�%�(K/x(�:���Hy%�a��g"�B/><�+���s�L��I�)���=~ꑸ(�����4����/��7 ��Bt���3��f��2�?�0����^�m����ME	��ٿ�˰�OƟ���n����n�r����l�@T���M:�����q��J�����,FP�9^�(��4�F�I�ǋG\�{�ā������8�`4�� C�o�s�������Sz8����1�=����,ķܲ�>fz3De	�'8�:H��#Hg|�)LI��Q.ٲ���������������_Y#�F��R�^�Z�� �[!�'���O�x�3[�z�2.o�Ӭ�j��x��H��p+��2�TX�H�j`� "D�`L�Η5]���#������PŨ%�Vo?{�+X�N�]/\n{j1�:��6yEb��wA��4PCYSvĐ!!ڎ��)X��8]���M�S������p쭘V�ZP>�
��3nt�j��'6�	����@Z��#Qt��7=)g��!��.I,>x�o������G�*q�-���rZ��5�����Og�K�=��u� �)T�]�q$F�u�������O��iU���S�Y�I�M3l�~u����@i��sY�?���eA��Eʝxv�_տ�
s5��˄	�`&�Y�&���Y/���丒���=]M��z�6j1�gm�Q,� .Uߦ��4]�p�\�!6E���fWL	Է9��񓯭�sLq`E��hʶ��?�V8�BV��!eFg��.�������~��`f���gYuq��i�Prb�os��x9���C�C���U�I���W�s5�OEd��b��od�$|��44�=_Ꭽ``����cN�
rr7:�e9���G��;��:��׊*��_ӡ��Qz�7�r��1�0��9�	.-3�B��~|�	���hS��&,p�L��-�#=�`[��f2��h`Q�q���a��d" ��#�����_�_�d7SZR�1���.K�E�A�yi]M)���(���r9�jd�G�V*50�wɹd�[7���%����zsw�
D0��/X��}�7�3:��\��UP������95���Q�����͚Z�C�̎�z䧽/n7V���A8���\1��I��0arӺB^k�����r��0G��R/jal?(Ǚ���l_h�H��dk5*�B���I:�D��c�����c��Z<ʃ�\E�@�b�}�j�5�tc ݂�aVj��j�������9�j�e0�-^�  �]rBU�&���'|<���G���k�PO�5S�����CF���[�i��o���*�S ��u ���H�i|���/�[��&�w_{�l��SjfR)"�#� �����L�z+�n�|y!$�W:�
!��
qa7�[�w�� s�8��ړY��t�k�ǻ^YĊ���\�S��?���_w�x�P�".7�E�z����]sL� ��8i�y�{��d�:�*���s��"Sj�U=�p´�PM�UO윮�K��}3����	��n��G�Zy��i�ﻬ�ٕly����E�<���?.�-�6�N�E��"$�<T��d��t�Qp'��G����4���5�C�u(g�]�>�9l���z��盱Jz�I :�#������O�b4��F��'��Ǯ��!	ͺ&�L����r�,gһ%�	d��e��(2�0�Ӂ޸�k�G���Ps� �#��x����P������qGᄌ��Q�p����:IĎq�L�_�^���s{A�L\z�.������v�.r �ֻ����@3�J�?M$�bzl,�$����T?�;��@�b0��� �D�x��3��L˸�O,fV�����%�>>3��\�Ի�9*/�\H���{�*I�iY�a)����d�|�²Yl\d��Y\72��x�	U	t.�(�C�hc9��R �ܚ��2�q$��@9uv�.����y�,�O'_��"�g�8�[�u�]�8Bl���z��o��,�����c~�p�(��Ia7%B��f���c�d#�,�%_[�`yT���|'G���߮��9aYf���uұ�$��_����E�C��f�rH̞?�5���B�D����v�����^}��)��Q�g��նO�D��QX�w�qeX$x3�[Qq�)n��	�.8���T�ܮ��!�7�-��ŀ�x�Y���Jq�Ćudƭ�5��ƴo_ ���9�&�W"y���>� o�����9�2g;(Y=�-r5�`�,2���'�*El"%��5C���V����mT�a�;��e4E�J��Z���G��m@���>ͅ�t}*K��L��Y�TCkTOlm}����t�Z�E�_<:8W��{��|�/,�����Wn�����L�����z`�<A��4�gC����l�
U�ix��Tӿu�Ї��ZN��^n`*��$c�w0�=���aQr{Xɤf^���0��Q��4H�X���}|�tK�qdR���Х�<��D����(�r'?��6�=�r�����U2/(QNH)TJ\� �|��Y����ō�М�&4�B7^��Z�qQ|�A��=r�e��¸� Kc����͛:���h����e�������8�� A�S3�z��+�k�?k�/�.��&�c٫]��w_X�*Q�F�b��Zf�U��2��Ȝ�p�\���MxH�%v��Š���K!����OGO����C$��y�^ݗ���cs�����:_V"���v'	(ڵ�q��}��C���lX�,��˄�Ƿ���QP�%D9{ Q��U:�r� |�e��j�iq�t��iBs7N��cu��)��ns�C5��;h^���PR���Nh�����T$��rV��;��+���*�i蟅F���:��5PR��[�olA����)��#`C(H��$��k�c"L�Zaz����.���3��:Z��d��?�v����Y�_���T�eUJwZ�B��6������l����������D*0���]7�~Ȣ-�<��n3��sa��[D�[v���<��s0��C��*CY�$�G�ex�ށ�t��X�}$?TUN��n���s���g��쳁y���Ya
@��M5��y��±G��������. �4�!�c2f��%�:�h���"l���������;1vq�=2�ŝ�B���`'��e��ڸ�v��y���ښ*yY]�`U�u=��a��t�hD���?���ʃ�P7F�>\k
�wt��CvB�5UoM1<&,�L�]�����`�l%�D18��C�������D�C�B	��4�M�	=�(������XW�~��?�T���9a�`jk ��q���x�r��� CݰzϪ��FF�0���f�e�(c�)'�w�����	6�c��jM)��ٕ����O����ƍg��z�3/w���̻�����ϖ�5�l�fQ_�WI�0v�]��p�GQ�|=>�*��Ga�P�r�S;��~ �2����g2,��	Ev��)�]t�Ѓ�/����o/�7?T�G����o"��M�}CB��c
0���2K�	� ,��8�[�q�i[޲�g�k�Q�����ڄǢ��]{v �RQ�*��D'7a�2��eqe���ִm&�� �sϥW�+Y*�d�������1�d� �m���Un� ��^ּ�~�ֶ�{+Ci�L��'-���9ث,�����Y�%����Hfw�LW���2�Z�bE����IѠl���3w��i�c��I^zv����l��n�Urok-���a@�����L��6ᝨ��#;x����R�;�E˙z!��Ϯ�ҩer�F�-Yn{ڸ���=����@>!ZN��K��{r�<�k�Ut���j��:�r���Q�v�+_���%�7Fc�ɲ�U2���������v"����U 7�C�u��܏c�x��}
Y<�������@D��ʫ��O	2�6� ������(��'�/oZ��p�(�5x�*���m��Y�"o� uD��{�&����΄Ku��b	��Ă�[.ԫq�yd�d!����Sb�������9��Ͻ}ea��e��Ȓ#��+��[�����d
��!.m.���g��"D�D��@q+h�$�NU�Nh�����h=NL�ƃ�����	�!HH���m�4��Ȇ4Oo�NɟA�ss0�Cv����H��!M�0]�`�>�	���(Qytu\�Am>;�L��������d�"T��
C3Ӹ��r� ���,rd/	���-W��$���2�J,}�|2H����HI�!<cI��j��ug��x�m���>��؟�x�:�>37���8��0b�;�{ ����*!X&l9��,���N�����`H��U &�ч������tj�����`P�i�Cg(\l�E�w�<`m�����U?
���Í��Y
[��"���	�����J�8�Br��AP��c�2j,n�Qp�˛S�]���2����,�?x	�����g��X��0_�M>�E�?Oy�c���6t�-:휧�������p�f��	���זH�˽�׷�IE���3d%K���1g���c��oRqMVm�v4 ��>� ���)L�g�	z����nd��,�W�������s����sH5o�,���b�cSi�8�\^���:�.a��{����'�Y��R�o�9��@���Jv�̿1����K��ؙ�%j!�)�~-]XJ����ĥ����K�;h�y�>�Dq��޸"VS=�h�!��b�
�C,ef�6K9���7"�XE�ک9W�yΥ��ґ'��y90F�#{�J�
���tbj��D��6�󑀏� �w{}�5n�����������^2r�V �R�H��6�"�%Nm��{ƛc� ZK�5T��-�q<��)q
I쬍TA�!L<���K�n��?��b�r��#>0W~]$��H ���bG���e۞u?K׌�
��r����)������(5ǂwK�T5E�����S\Ϩ4�7i��u~JI���ڤ�?�or!۬����af�U�
��NzFצ����=?F����c�!<J{,��W���3���a�> b���KM�;�ΰ�hQ2hn�`�	�F�H���$����}^j����wn��$(�a������(gP1�ŝ[U"d�j��S�ǌ� ����99�.Տ����Z��8�=@1g+P7E�¿��&V�v*KPZ%��Q�t�͌I�2V�āzGjy�\;����w&"��fp���'��@p�?nBS��?,Lg��mj�^Fʹ���������2�z5��
�-H�q�xX�z @�(L��+跺��.nI�����l��/zER2A�(�߹@�
�p'��*�yYn�H��C�긫����^蔍�8�R.�Nl5�ַ�S�����_�y�!y9A��,>�!]�6��e�\H|����,�om�t��ZOW��t5šN/�g��ᨃ[�����yb��rF��S�d���'����3d�B�A�8�������-�> X�s\N�Q�֏VH��Н�I�l]�6�
�Mn�_�A��\����I��:��6�bq� ^� N��e��ui�gX�#��D��8�V��3��ek�Za(k�h#I�;�����݆æKm��e?ضl�}�E»>�υ�B�^�?�O(T(/^���K���u�����g�3<S,�f^�ⷊ5bze�zt��l�`��Awo�7rF�Y�+�E:>��_�v�
:��%aM|�WQ�[�n�b���G�������b]�R�Gނ\�uo�4�&�����m��x�煘��	Y7W.o�c�j��e��nI�[l�I[U
j8ц���0l��/dr��5;j�h�ð���ң�9��D���c�)����/ j2���TuI�d��gn�S�]��[�5Zfq�/��
�2#d�0�����>��B=��$6X:��h/��{ag']h�D�g	�#��2��Y��c��t��H�^�"J9��U3�9�]ĝ��M����PC���"�d�!�vd�>5E�=Q	� ���$�2�$� [P�Z��֡�2��b��V+�C�n
xއ�_�P�[[Z��'L1t���W8ĵ3]T�C�-a#~+�Ͳgmo\.��,����c����2��g�P��<j�Ss�d����
7�C)����A��\t*Ǣ5]�Z暚�Q��Ov�
�d$���-�L�q;�U%͵f�4�n�i�ߨ�G��~R�E��Pb{�u�U��?�Y�c�N�j��U:H��!��]�9�(��N<P0g�`�s���f�Ҿ��\��*®j����l�2���k��|�m����.'�	�5�N�ey��%�6�)6��ja(�gU���Ǽ�
4�m;�n�q@.h��ON��j�)Ca�����0sV��U��X�qL?c��9���P./�J>��@^�q�
�?;����G���DW!S��(�V��=���J�p��-�4�� G50̢�ь/���P�AcW��@�y��>�XoT��=�݌��~A_�	A���}^�Β�cy%��B�`�k W�OU�lWa���楦����'��\	���`�䖞�gb{[٤l%�����g���+|L	��7�h���x��޼c���RkJ��v�4g�QqςX�i��A�t$��]�kgg�/���EP
�Ċ	#�#1�J}�F��j����D+��n����8(�\	�$�k�?�#�4]�[E.�=���É�u��ȣǵ��LA"������P�8��@���}\Mb��i�=7�Y�&�d zR�-�'�C9�Y�R����j�x�f M�>C''C��!�� �r�xG�4��uFNxg9&�'�ܜ�{4� c�������7�؆`W�@���.�{��M�4-p���&�2n�rK<��l��&@�F(��s�*�J�������e���)�J���b<!鉬��˞l�8��L�����8p��q�\���qT׷��N�[j�n��l�$w<jά����Uo���:�b.Q[Om�z���I�Z�&��O^(���u�V�%����Т��[l_8+O�'e��=+��b��Ĭ^��ۧc5'��5����_�r]Q�����9���c)6u=GQ���	x��\X��L5&He|G���/S0�dY��s�_����| R�"6#���V�ӏ�/zEgKү����g@ft�<_���DfZ��+����8�0��C��l����?"�VPJ���ü���a����h��P�A��rö�\��R�9�󍀩���b2��E�y|�m��,�@ژ�cb�gTg�K4,�����@�Y�[�\;�S2��jJx?+kt�S����S��M"!��X5�Ʒh�],{7���`��#��ך:�˼��~�������;X�yh�M�u ��}+*����)@duA)i�Z��)b��Q�v�� ���aCx\��$�b�
��C���t�2�dDfE�>e��g��������:�Y I�E�HKHs��,����Ds��[��+�žoK�d&�.��K���w�I '1kw<@�`��n@�yE6"��>!n��e2I�C�ѫ ��իͨ1��p��W"g?n�������o}�zO;O<^���/L�GT8�OF�P8H	�G�����fƄ���J	�\�.������{� ��@>#�a��l{���R5'�uX�x-Wv���VBIz��Ͱ��˃j��;Y��T�Y�
�X���Y�h<�76;v�fOx$�h�J�j\§�p�������E�F?��9��8�����,���J7�dNy�pL!k,L)gI������S[�m����2�p��T[[r�^�D��fIg��2��|q��+��gt�U[�*j��`k�#z�z�\W��z��59v*d��L?�@'+p��d��$���r��^ ��(IJ�����]����O����m�`a␅�>&�k��JTr����-�Vwn��u��&N�~eTi/_%�&�vF�������@G3@�����A���؜Ʃ�	���gL"H�ƀ�e��,��ρں��a�$�5�5G�f ��b97/{Ώb�7��*�Lj���:T�m��Z��������)���i�S�F����x�~/�1X���ƺ�PJ��� ���I��BP�d����S�������Z&�O`�7��$ߍ�
X��ft���Ni��*Jxs�+4�>ߞ��]�KN�r�A��M�w�"� B��kCq�hoO���ZHg��	/��f,.W
�2�Ub?u룰K��=�v��2��sZc��$E��������[QG��+~�ec�8r	5������K� �ʇ�lk%��
�{�xP�B��"g,#ܴF���{�9%:<�{�R�9�?����W�JlϘ�d�H�'a����j�|^�M_+�M�xȠ�^j��m*m������~��v8�'�,�%'�bǁo�j�:m�;M��BD�D���3��v8�	�
��������C9���r���$+��0l����`Q�J��'C
�*PM�2�ռ�>����"�-LA�c�ݗ�C��tXG�#R*�p>�2�1���������x9�����8�7P���q�=���YD���H����$��37��O7L3H|��������H�YLuq�����k����|��n�ݫ��e"�zO���<s�Դ�fS8����D9*�'��8��!�SsŹ�eO�gl�dvC٬��*Q�~�7�T0�0Zu?־R��H���#���̦P�q(:r,�� 2��.bs����G�zt�R|�v���-d�;���5,{�! QHZ*"NV�m������:��TeM��$�C�2���0����N�@�D�G�f�o������|~�^H�;3Ȋ币�[�?6��z#���G.KV����U����!r�/\[�b"��`�f�s.!���ܬ|~�-5'�^�^'���z>7�'}�*�y��U���r$߅mvd�ԅ54%�Ӽ���נ��	_�f���嘔���2�0l���ՠx�[^q��ӂ�l�gv%i K?ޛ����Rw5�f��K�Ⓛ��(�Ɗ!-���g7S�`�8R6�E�p�͒]g4�HTہL�<�KZ�!���o�Y޿�$&?��vy�y58��'�t�h
Nph�qQ�,Gp�yx.�(����B�Gۂ��K�Ԗu�G[a+���wl�����`��p-W�ca������^���T1���P�b6���؝+��'4�X��B:�"Ʉ���[+U�L/�n4��=H�<�8�:],uw��-���oG�>��3�g�s;�K�]��fF�R
4m2�KHh�x�Y�.�[*t:YK��- ���o	km�Y����{�0��i���4hp$O�J�m�6#��S�7�b��"H�A���v+� 32��I����i����p�O�)���=}5�C�#�F5�W��_��F�����Mi�GCB�>u����YXL�y���025�M��C�.`�����s-21F����mT�g~��;��Z7A֑�9t���.��N�\�IƱ;m*5*W��,��'*��G�;際�CR�q5s4�	����A䟯�I4�N���o���]���ڟa�P�ܚ���t���c���XN�.���\�t�e�X�g����b�b�����ȵ�?��Oj�Рn�����?���xW��w�v�e�T�2E�2��X0�i��.��J.���u$MznӮ��!U'Ȼ�Sw�	h,���?�v� ���F�y����#����3��д��p</��Q�@f9$�:՘H��
���z?�3I��zT�@`s�˂��.�wJ���;����8�M1� m��1q�L�qq�&��;.u��q ���eF{�nwYH�����^�[��z�$�<��3�����ny���c���I�q���'����^y;�R|��ˡ�����i��8��'缭����4�����})���wnvNcQEz2+�a�3'��@`pD*`�i�F�Y�,%&Ѓ��u�� MRnB��~G�������2����s=:��)�rK�ӒV��y��
����V��x7d̪k�Q�u	`�v͇@�Կ�
2�zwf�C"��;�����s� S�,M�x�l+o�"q�{
 ��ևs2��"q�h���%[�3.y*�M6�q��Z�E:,g�5N-i��4�f���k����`���Q�0R��R�w�f��h���E���ǉ�e�TE�E�<0�^�97?)=5��ZAݹ/���/_7�T�-�Z�L��j*�G�\ND>�`�U��^�@�	e��*r�Ο��Z�Yy�����;���ImtK�N1�� ����񩠬�e$C��#�d�zߕ�3�kر6�#m��Ӄ����oo�0�jw`ʧ��s��N	��N�C��ʂa��X�4�(��!�K���Q�<t ��Tt��a%����b�������*@�"�E�W4/�O�x�庴�����&�(�O`��rԋ�e���/=�nr�%�0Y���ڭ5Y59��#z�R��K��h���6���������6��Ͳ�t��VT���*q�2OtsÇ'���Rꁗ4.�0b��1]�(��_Y�5&���� �ϒdNPǨ#���*ċJ�y_{^�cH��Ee�L�n�����,9QxZ��Y4��GT��Q7��Qb�)v:TB��m�Éi�?��Z�,�l�~S�зY3���s����K#X�8��\�f­/s��p�c?��U�`��W��'�����
�'�W�z�<(?�	FR�e�����c�Z��RD����1��tcñ,��)i�y�=��̦mk�l��?����Z��s��sS��Y?9��Au�=�X�������y� {���ʋ'�0f�DM�oh-=�Sec]]a+����D� ������[�:p� Ü��{��K��hJsfD�v�0O���K�%��?B�oc�~��!Ip|���-�U'��B$��v��x�=�P��B��m�����/n¸VR;���J�))�U��{l���ɷ�}=-��5�B�465$�/��"䖪 0!��f[�s��pY�b�O�/�6�nr�
��G8R�y�+e�?x�6zmѳ��e|���Y�Z�K�X���
�M8�t ��H/l�g��la,ʬ'}�uMh�(j�0��)h��Lw7H��GK���g��я|�:���q�a�8�Ÿ�b��X#B�S�0�m����p,))�~�M�xID-t8Q/Mp��#{�yTEQ:u*ܯ%5�Ӵ^�Y��HOn��Mz� {W��x?a�sgS������x���(�IҴ��x�+	+��;�c�j�׽Oہ�d ����x�z&a�aɦ�ծp�~lϺ1��9���bz� 2Cg��?gA���$"��1�`�.<8�68��̒x*�Q%z!&��L�(�����o	1p���:�{����g-���Ocˡ��<"R���ָOؾ�(��z~[�^vM�V5���.@G�!���L��<P�&�Hm��y'���GQ���.~��
`R�	<�m����iJ[�'^.y̬A+F�fa��n4���w���G���B���G�(�a��^y��o
Ш��"�6�R�.����f����2INkE)�/��m�8����P� ��v�z�D
ʶ��h)Tm�-�=X��s0"ẅ������rМ'o����,����6�/���%y3��K!w�
�I3��\l�P-��"�cv����S�rkV���L�[A�e]l�G��3����]�8��Y�h�F`�aI� �����1�!	k���r1Ck�l�2��C�vr��9�a�S��ԡf�&�;x|oф� ��o��(�;�ı�H�6h�#�>�B��~����<���݌u�>��V���tuXd{8#���R<C�칹����}DGM������P�W�^�J8ft�N��ς���*�l��u�te|π�v ��đ���Y��� 	���c�+<H�`l��&#x��oM���\a:��5\x� ��Q_�����������LN�o�
�	�5,�1>��LS�A`��u��; |�Dz�{$`�7�L;/�*�;ʻy�$�{�O�I��m�����~&�*�+��]���s���5�?ﱶ*�s�YRx�֍��K ��'^�ຌP���#���϶�iȝϧK��m;t�4�oY��L��0��(�-�����1�����6Oy��6P2�w��y+�<	�L��{�7�^�bk�O����>}��)�nE�"�^�	��RI��騞軆��ڥ�43p9�!��'�hz�νo�w������Q�1U�`�2/b���t �,pwv�@��V�p"�2�r֓���W��<��>��o��mAۺ�;G�P��{�Pzi��Ǭ���qW�
$C���.�[�4>C&�9!xoj�,�Dav�"BU��nJ�{x�Al~�[�	�u�G�� �M��p���F�I��w�V�8�]V��!�j����w�g�.1B�`�;jx�E��ElZ���������C噠�.0��r��@���	�I���<�n��#��=�0�ؑ��wpj��vTw��X���:L!8׽F��QG�
n�3��E	T�ʹ1��a�������5�+���}����h{��U�7�m�ieb�@�r�%	)���s
���j����1�-l�v�=��ys�C���#u�
���/��9i��>��)3z�eB�&U[��²C8�x]c:�f��Ծ�F�	���B��U�pg�t&���u�:L����av3v2���yY⨍�麏MP���J�f��
g��Y���OX��ն7f�F��:��	�7�T9���'^�S��<S_Q�c��Rav�迦�h�o���Y]/�G8�N�i��&m�!L�O_wL�Ȉg���|��Ś�I-�GgҮ�,���GH1��Ϋ�5�T�tWU4��	�*6�C�]��}M5��N�=wL���H���%bގm�12Gn��[W��vt����2�pr�?���h���]��Rᴵ��䟌$�i��P��}��J�B��s�D�UL��`�����]�+�$��	���?�]�-��,jT*��;�^��JD���5�G��Gf� P�� Z�|�
��#���$F$R4��rQJ����8�Yd�_��[�}<d)[���b���teL���p�����ր�f�1P���5F#"��cSJl�Hd��yKpo*E �G;5�`� ��#�be�Xb�u�* b�|�٭�>[@õ���)��?��Q�<s��(F�W��d���5��Ω�~��BS����-�3��mi�.����(��~g<����.�,��>8I������ܶ���!N A/�_^xD�� !�	D��,���k_$ʁ�y���YC��;�
2�ρe��Ps@�����^��n��<���z����p7 �V����:=�,��6��_�Tt %�SKPkNҠ�;S���i���H��]�5�}�A����隰��b���@1��W���e���ucW�,RaI8g͓$x�%�E����M���GŅ�L�mӣB���^�L��+��t�?��G��Yȴ��Q
�6�7��ïpmZ��0oDyj�ODif��O$�b��Rϟfz�~EG�C��'�ނ�A����/H��I�/�g`A��t�b�^yt��,���xPs�� w�~�m���UkV�I��<HmԄ[.x��!,cc���rp��UE0����#�2���IVP�<�w��qi�]�͛77)����C�/,�$j��Sfc���b| qd�0^���6�����/�Z�=�^iM/�YU% K.���Ic���;�?��ap,��)x�,s����;݇/�P.m:$(+�R�ʼ�C]"H�b�PȎ�v�́f|s��F3�QIܘ$v��D��o�a���q���p%��@Sfz��GHg���d��kH����H�8b���� m���\�w�u��J�jf�
/���ʉ����K�c�B�˼j��O��|rg�� kIi��<l���]?����Z�t�`�[�������E�ֈ��U}�D7/����#h���0S�e��v}?��58�	�G��[��Բ��#�7�i���Cw��sC;҂����.hř(�8����h/��g�Ӎf����x�������$���<��G���³���R�CX85��L5�k��y���E.�L���&f�/�t5nvWjlK�A8'W� ��G_=�b�h:��'���7`A?c�c���j�f6���v@��Q�K�����m���<¼9
'��^9�k�*nztd�����	�9��Hfsǜ���%�����̾9�_�	��j"^��>���-��j�x�54>�z�����s�-�4���G�jZ��{��V٣�g��`�	�Ł&11��0xUv5�fn������[a��� �}��pl��u�f
;do��:|<�M�y���u��äz"���ދ>��K��փ���ҭs�b����h���HEBk�r���8��L�矼f�̋C��@�����?F����Q{{ Fө�Gۜ��\0�����'>�M%>	�; c6�'c/Lv�'�l�K���q���\����4z^9�1�"n�C��|�̱�:C-��x�b��Z|Y���4J��V>�S(�i�4�0/_&­y�6ٿU��Di�ǆ��n>��v�?�&lXq�G �L��������nXP�o득fum�i
;����W,��7'ACCC�WҊ��Ar���=�n?�.��ar�[�3�)�uI���xS!MU��͏p����!DLRou��h~��Q�
m��i����du�K�*b�{e�H�E?�AW���,I�R�M=��ߒy�iՑt}G��L�C�'��Z_�yG�%8XgYD�q�c����?�:q	#��zޘ����z�:T"s�B:�L=2}{� z}��*�WN���.>~�T�ه�ɵ�B���/:���W����'j"�'r{�\��';�Oa����[����ӤXL��^������zf .�r�X��;E�	�-k�e�JΡ������,c���Kni�d���a�G+`���!��)+7y Ӹ�G�DtN.�h�<e}5�h0�ꕧ�9�4Ϡz��	�_�@���'�?�('�L�b�YG�7�O�p2
��A�C��HQMl�O�wS���<�:�9��[fV��7>��P�|��������w�o�%�4N��I*�s����S��˚fd*+ >h;�a�r �3L�q�uX�"ɭnI(K�Ao@'��rʏ��^sy��!���N�9� �1R����ÛHi;���{"t$���%P�u(���6�ۖ�JE��Ϊi�ڄ'���D"�\+�J␪��<�𑼟���c�|r��͏AR@|v1�Vq��ۘ�<
f�>Γ.�4��^F^������;����>���U���t�&��ӹ� �~�8`h���}�ݭI��[wO�Y.Օy�Z�26�I����h|�2z夞C���URB�f d�b-�����������9�x�X{�,cQ�Q%{2JAӵ��A'��d>�:�uس�B_��K�í�9�̋ p-�J�F�j���:wq�)hn"ug�J#�	p�}8���eo��$�<m��|�l+W��q�i?��r�ǅ��wѳ`���T4�Ʃ#�t?�,��4�ݏH7��I>7�@�5��\���Ơ�L���nhrC��d��������$0>$�\[�ҳ��j�|��iV�8	K�k���="���L�,���ߪ�g���ZAHi��fƑ�����QA��u�7���d	.{�d�<�P �(z��AX�ꚠW�t��m���ʧ��>̧S�%˾����!��冂�S�r��Y�Q�^�=�ʰYtb��������3]H���% �3�~���������x�r�3�I����?3���{O�Y�ByF��%�~"�x��s�o���d��茖Q���5r���p��x�I�j���!)�*��_�:P�( �m�J:�a��B�ʑ�1H{P/��:/~:����c[�s��2e^��������x[#��G������8Z�W�)��r|[KgV���QK�#��6n�{�I��b6�g�a�!���p�^����j�OPl�I���+5���J �*���b���}G�虏�&"���~r��xj�A��'�D�VD9�#���[��d��r���<׏X�|�;=��*���%If@����޻��1�0b�R��&�E|��>�4�ٻ�nS�t� $">���hF��Y8ls���'=r����2���I��h��gEZ/���׸�o���BG��S��g���Mi��ʔ����]`Ƿ'1݌쥹�\��6�7D���3H��Yז�^��#��+3ZA<p"�-�'1����¿��A�H��+0�sj�%�"�+O>��>�4�0����W	 SГRc+�v�>���ѤZD��7��~£����˽bF����=��X1k�����p5ޘ�Z5��w��������}4#2�՛�9��!v�HGͥ�Tl�|m�jڪ@�*�nx(�^���f`�
� %]WUzi�'n[�<UvA~��Q���5�'���G��J�D���$N��C?K�r�c&7����~�-���Q�����A�=B���D��8[�w��'����<�!�J�1�{lkY�?�4�$�j�����\^�����+R^im�E%�<�����~-��֧^%������b���+bG I�۩�%u�4������i���w��ln�_e���������-ew�9��d8��P�_a9�Ǌ�xeqv֢IPW�"$2���S't�i�`e���F|�i�{�X�TiV萎��"#��	�e�������GZc�v�t��|:�)ٽ��5ׄ2�84>�>J�|Z��&����ׂ����SM���j��[t�|��3&�1*�������E�	9�8�m�,m$�8����]#������-���|�&�7���P<�#�{Mv+���(|���'~�� c۶L�Ow�ni��#��k��ni2qn
r_�I��s�;�&%�YǪ��\}�q��4-�o�>�#f��J�K���;�7\��U�Ɛ�f�;f$�^c�a��h�㎄\v�>�a�,ۮp
�������$����>��sQר ܒ������rg��#[�B�� �Tk�9��m�Uߖ
	�iO�*[�.1��6J��˻0�}�ƅ�b��!>V���Y��S_þ�I]Z������k�|��>%����䀞��L&"�&Ã!��"U<�l��哏(�'=�Q���BZ��̢�Cf��j��uí�qW�]ʌ��.�L̃��8(���[�4�� �[H�Hic���Qċ埔L���|�jR���D>v6�$ИSO�	'G�r��+W�*qZG$/���&�0�j����T��:J�	�U'Q��дٞ�[&V26%�*>BF.?L��� ��kB�+ʆai�����V�����k��k�Z��'e�"��cz��/|�N���iٺ8�ϒ��(��:�Ab�v��]�Pzw{N�ġ�O�&z'ϵ�|�QxsH�]C���"2����o;��G��h�N�B�cש;ٻ&!M�'�Y���6m�֎��(�
��� �$þ�Z 9��p?�v}��N%��%�J��H���]o���OԶ&��[�^��,}��ٳ�m�|�PZ|��'���r	o9"�S(�Sb�#WK��B���
�,�ҕrW|��j&�Vh-�!��`���1�iѼ�Ei�^�S'����%�A�Kk>04��ӔW���$�,En�gΣ�����u���I5���9�Sa���}�ئ/�֎s���%5��������>W$�ję*�C��AsVN[zݢ�V'O׉���K'��t�^����[Q�]z����a߆��W��밄���|��垳�
e�EWos��^�B�A�{�CAm�"�x$���X�#�_<Ls?��03S��B)���8�V3�d{���Rd��+3���"~����ذk��,�����i^\�����m>���]t����C�\x."	a���C�
rCkf�3��Ìg��</�31U��~����鵦�8dp[~TBN�3r�Vٯ�[�*�(��Lx�"��f�ƽ�e��Z�(�E��$z�`��$gY��Ɛ�pTG{&�ϑ�(��p$a�C!�.�]��(��
c�D`s-��b@|���?�K�jk�	?��7���!���/���!���ù�B�V��.��=�zj�:ķ�y�9H���>�&T�b�[�;\3��}ƒi���RJA�}Np�{㲃O�>����E���6r/� �VE����]y_D��l�Jϥ��sJ��r�5��ART�o����qǰ��+F1��2M�+@�p�U�Utt�@��à��f&�ɭ�;�yh-��zѿ��le�4��,��O�?P_�4��AI鼁s� O(��.��g-�6�JU��Z�W	�x�t�.2z�mrs�)T�ƌQg����Fe�y(�<�o�P��~j�6�Z��2��%�?��̓�r��a�����p�6�׏��J�`��AN{�ui �-�܅=�
j���xe�&�L�+,#:J)��ψ��=wp��K�+�u�nƩ���"�h�Հ9eEǮ�PQI�u�[\ӿi�]06h<�F����A7�7O�O�~������-�|ؔ�Y �=�A�#�m��q���;��_G����fJbԦǙ����Ӷ=9o⅚hyZ�xw�.AQ�*���@�j�^_���YO?��|���.����+@w!ky����Z�-P^�+<�H/D���Ay�BZhdJ�o�����*�N��*�hs�
�,PX[$(���"D�t_Qt��o�����.ѯR97���#]&r���O�&NK�<꣫2CRQ`V<���//�izn�7�O��O���~�h�4<ї��ƒ�>K�>kM��y��m�s��AN�0|�;>�@&���(���=�B�۱s�񬇇���y
J�o���}]��u|�3L$<�Z	B*C��VW��@�C���J��U6���ѓ鈐:C�Mh"5�~������5X��wj`f�^�����r�r�9�����k>F%��>�PttN��"���>Q�c���YQ<5���7Z����oF���OX�E�C���:Z7r'�Nm����061	�nf�{�tl|S;�6"����\�ܮla��H�{�>����ɢZ��y��ĳ, �����O(����W��[�JD�t�L7�O��Ng7o�I����9@[SZ���)6��N��X����}�y�����elcZ`�$T-�){!}"��wzdֵ��7y6ڡ��(��a���퍕�� 򳐢I@r;"��1"��Zc���ܛx��+��7�W���\�dk�w#���n0���Urn7?�n����`�<}�l��M%����B'����`8pRX�� � ��5���D���H4 ~�4��b�s�C�m�_����T�E���HW��E����
xP��{�Τ����.!�S�XK-~��	u�r�f��i�����| �H���(ۧ�sz&�!�RAP��F�.A;���q��%Ri��;���U3��jSt�+:Yt��n]e`$v�,J��c�~w�V�B�TJ��@�1�t%b�H�S��!Ce7�K��~�e���#���o��'�עNؘ0��a-��;�E��� ��O��{bSovH����/�{���ˡ��]�Jp�~L+N�Yn1�������`(� e_x�<��}?H$gK��YBK;�=�����;BП}��}��&�Л�=�fY�����{l�����$87�Th�&>�q�۞�.o�ā&�
�+�-S��;�XRk�����|)^�@�gR1��W/��A+�T`���Ab�.s�P�,�Dm�rK
�k܍(<FG���8����m��+f"��J���CW(�&��v��j�,��Evy��asޜ����`����*)���]����f|=��V7Qm*�6B�6U~�rf�s�O	�
#2~��1m��&*CP2�M�X��@U�su;���Yj*l�T|�x�SZ��Yת�E 
{i%_\ђ���V�E�"/���=��B?�¾8E"���Qs�K[#;A>��{�1N�/�����ƃ�e��lyq�����p<�����R�B��F*�
<# PH̦��6~X����F ��*9̃-ދ��ی��Op�L��o��� u��֑�e��hXe��<Y8�_�1�V��b�)�;Z״h��ج��� �l :���o[����y(��D�q"�w�8%�o[�҉��bjd�j�Ŝ�*�����<� 	����#�.��!�����K���a�O�lD����/�4@��&%�*��!�P����POIwq^�9
�Ngrx��d">0��u@H���>��QATN��Ci���b�0Y��,7��U��t�V�80v��CsM��U]!u<2g΍\�����	C��7b���=���S�clrl&�> �"O��a>$l(��v�N��u��h���%��ь����JD���r���j!i����6���>�-�:�r4=!.� ͬ�i�0��Q[xC���Mwtעl�}W^^�f��L�����}N���)��8����d��O��o�)�F>�k�c�6ꁕ�@�Dd��w���]�&�B�K2�=�ʓbQ�0�+FU��-�m�Y�D�t̒Y�ה>R?"�-k"�CS&y�b��a0��(�gf��N�.��S�;"�֋�b�������\�c���HԢ�o`gw�l9��]�X{�m�ߥ����Yg&g�&Z��,]۱GTxr`���qJX�Ud�T(�����b����I�07a��֪r��Z *��ea�$�����������h�����玒@0�~S�~<u�j�`M�EDgf�w� �I���T;W>ݘ�����uBF?3���1�⛦��6`�y8j�
ǽ�z�* �۶m7����M�~�
�B
^�"�"��}极- z>i�qs���>v\����-�Z�L~I��&��=�Z���N=�j�7���E?�}Cˆ�J~&Ͽ�����yϦ�@�*�Q�%p�X����e��G�t
Z�3�n�*�	c��J�� �ZQu��������NLP8���Oa�U��,y�fi�o�,����o��q���̹q"$Pi���u9���8�����c�M�V4�=iB��!��?,S�B���IFs�J�Hػl�"R�����c�8�,m��/Λ�ĵwuM��m��F��j<�$�И��w\*�����&r��UG«=
��
P'������҆~�O yx IT?��;���*�9�^�I����58+3�6�F���W%MsmN��2(lex�mb��;�����V����u�pܴ<��?����Z .��/�#3O�
�FI�x��=�h-��q�w���!�϶YLR���x����"jʻ$��NX�D�o*�췳�����0#��RWj��\G9K��w�Z�z^8R�5���ޚ����$/�q�������zM_^�L�#z������&ßX��Оg���[�	���˩��|��(���:7�7%�����Z/�����@d�y�eim�(���+ldynx@J�Z(6��oV�Pݦ�����]V��lK*�J�����x)��Gb� h�=�ّ��UmTTb&(�����ړ��������]��Q^����p�6��>��B��T'��ٓ�,��O��(Ki&�C��Y�b�UDH	�5W��0��SR�<�\�Ѓ"���3f�h�C怄�,l?]�|�l����k�,�HEv�A�u��o?�7�������v��f�(�� 	��I���'�/N�Ć�X��0���Ej�q:c��*b�afz��m|�̀�g��ѯ���ɀ-`�x^��̘y)a�׎�a��:RmY��6���.���JK�r�AR��������L��ُJ�H��lp��2�"����������1���Q��x�t�cģ`Z�;��dq��ъ���%�Y���rl�L����I�Պp\1f��#���!�hc��ӹ�Խ�>vg9-��U��9�==��G4���$�����о�I�YꜪ1ϊ,��O�QX���@���|�v�S-7kJ}�K�r���h�9�Y~y�rA��eU�T1���q��*{��<�>e�>ˁls1W7}�S@<��X��-	��L�p���UO~������ �J�ޱ�1�%��ƉG2�����g�������%L�������1)�H���.*o8	U�﭅Ō��1��������+ofe�R��.��k�k,��{F|��j�B�B��b1XJ�����Ո7����Ԯ�e���]�����*JZ�z�X1������U�-��ȑ�E�I#�?�`��H�b�����K- �� ,ީkN�=��)I�I�����Qq �K7��g�i��)�����w˼W�ʧLc���`3^��mgld@���y!����ڰC՞�,T,�y�rP/h�=$�t�� *Gs��6���O0'I��8A|�	��V)�6G����Y����X��ڑ˼�y�h���;�$!9������z�7�أ	�*���8c��b�fp`�V�].47����X��D6?*�g�*gs�hu���B�&.���,/��{i"�;k��Z���у~<�~OO��E���i�Z��}I)n���8��c���!���"�4��O���+��t���`���w/��@*��j��)CWr=��[��/��Q�޻�iG%���˓�HE�j|Vv$��i9\*��/�$��'�2y�1g~��$}��x=	����/fP'�F���ox��k= ���׆�fy���N�'Oeӄb.䈠;��K;<��n�R�).���?7���G��2��%�sD�'Оy?!qF�FH��d��y��]�Y���Q9�z%��v\xJ�I�Ə5|�U&-���똕�֐�R�(�X��Sk��9��  �զ���Y��$ګyI�^[�@8�+�' �W-�1H"�c�g%$�\y!�ؑb�c�'�����}��#2Y�R�6k�1!}��<�H��tŋ������z�|�B�_�ɺu���|�֞ѰD�W,`p�}y�4=E����#އ��`Q;�L��ݘHnHfS;dw����G�ދc�rW�eQݖ���4�s���jL��dʏ�R.�ԝQv}�����G�i-�@#�tZw��b�e��z�u���'�`Z��LT���[�ɔ�u���J���yw�O�0��π��&K�*���<L��b��k�ږ�\0�jSa&3NJB�ro�9���d\܆����O�-Uv��xh��Z-p��c۞Ɉ{gw���ڽ���[8pm7�*��7��M�>@��QZ�*�N2	ߨ?���g���/�O���>|�LB"�lj�?�8������fdL*j�i�`���.�F��}���OP�x���OF�t����r�$Ԑ���J���!0�&��o�|[�<J�Ɋ�Z�"�ձ%%�&6��BOe�L
B�%C�y�6����̈́y�tm$B�e�y�By�Q
�7!��q�t+ЀK5ظ���s1�!t�G�Z��xLV�[�B����(�2#e;y��(Q�rK�L�^MPT�����vy�O��X\�t'kø�b�H���Gv��Qqgq�_�#�� �!5[�L
������������5�>t��Y���VB�����D{��u ����S��8����Iy6��� '���&
W���W�Ls�M�j�k�zW\G�)g����	�)���0W���J�L��v�e*_'���O��~\�{'�U����F\3��F����q`�K���#��0��@����:/h�#~�imsq��~�n��*�HW��XP��P��
�	Jh��m:@t8(f?�Y~�Y�Bp�𳚛������๸��2��;��n��S��	S�xm��|�a2�q�$��w�sl9E~�o)`5��ON]W��
9��nv�*�T)��F��0�e�#~���~�ȼ#�&!BZ�Gg�_�&� `�v�֊��	�.���.&�͋��b�c넲F|l[��Yu�O��4Y�-3�~�A�������r��:dZ�>?�q7����i$Ӿ��"_�y��$��-�?��M��;���RZ�L�さ�34+�8o��%j'�V�̎^��F�������<h0�85����*zK�R���z>>��i�^�f���e|�Ò����GP+!@S� |?�A!R��х�X�ٷ2W���
7������]7���_��ۣ#=���?�zl� ���s�X@s�J{��I���G�b4+a��IH��$S4�G��qy=��0��灁[I�d�ܫ�6����Y�8�!��:�=A�;����ns(K��Փ:#�������G;��RDT��A��3��,�A9��u�E��Aj[�`-A#u�].͞����s��ڠ���� �Ջ�v�:�[���5��P��{I�D��Je��;�A?œ�CHJC��%��Ǯh]��	2���[^ht������z�atu�-��]�` ���S��f]�8Z��DO~�(��OZ�c6x�Z�Tf��wF�O��WEG����34�
��G��*��j-R#*�HG�uԡ7(�� S ��� +���y1Z�Ũ�`��25$5��!��Z<�Ɠ8|�g���TU :hsC�6^,�w'q\�YBZ#�j=��zh2%]���w��8>@(�<(\x��#�|�U����qxY�JrIv����d̺nV��ի}�Ʌ*"��i̔۞�i�ּ!���P�yszd���j@�<���U5�:���E�1�O�i�ih���>v&{�2��r|{E����:m?&ŝ�� ���
3-Xc�8r
�����k������8L�S>� ���i!�a<�wPb�k�AQ��
N��	{ܛ߾���S����y��Ee�ӡ����v;?.��*1f���k��9��D�6LB�wE�y�׫��s�>́�y96�Q�pT�kX��[az)@�SXv���Y���?�n Y�&�>���!�UBQ�Nµ]k,���əu79e��o;Ur�(����!�TT�)�<'|%���2�����:�f�g����>����D��B	�K���[��ՎW������R�>�	�a@y5���G4���=��f��	�����6���	��|=R��a/׎;G�s�'eN�=<
�����Jw>-�A�η	�n���
��s8e[b�������L�zZ�R�B���	U��G��y���4���w���E�ei��#��f ��S��u*� �����KLDk$�~����#�7��엧�Xߧ~LV�����Ituk�wn����A4��7*��<$"U��@NX+��FR���0(�&w�]�o0����qv�Y�ð߉��<2���[{6�����se7�S��[A�xm��Ȥ2��)�NH�R��hZ�S���@m�8�4��}�7vZsz���~��d�^i(���Zo?�(�k���CK3Sfi@�0����<,����h�n֦��) �����^kq�#���2_�}�9�+MzT_w�`���{S��j�c�(�͌���șW\��+R�x<0���
�^D_�>�C�;��G�U:�8���=·L��)��������<�n�"�U�-ʹR��Y���,��"������z��|0Ix�5/Ӯ64E�S)8��-)����Lx-���W�@�d.����D�Kx���mω7yU����j�{���?ȹbp=6�1�e��%���g{�ŭS���j���Pq��IEhW�$i�Ʀ�z��
<�8��x+�Z|[2�׌��;9Tx�c>x
Xߦ�Y�h��
��\�����޼4��:�3=>�pv�O�wNo��
���Y&26����l%��:"�S�`�mO�$�q�[2Gl�h������'��{dyE ^CE�v�Q���D��z{��߈�us$E�3��'lC<�_3�E�'81���gq����q�0h�/-��he?鉠�Ai?���B4!�i��B$�{���R�B�B��z�y�)����q�CN����xlW�4�F��q_!�	��O��$i��C��:������-�߸���,7�E��ܡі7��&���p��T
�a���V-��.��9���@s��IQ���B��`[����[�Ww�Li�/�_�aG���9���|�-�v�F�M�?�On�}(D�/J�%m�]+��v��5C+K��]i �2��|�8���`Nax��!NPy��>��DvQ��m�J�}4�q$��Hp��[hSw�8X���w	�B�rc�w��>��_��y�Y�V��#`��R
���h@j\6��e'�Rb�1Z8�΃��7inp����n��]�.t�s1
8̞���U}�U��q��)v@I�4�dc��E
��9�����Cˬ�X{�^uN=^D��i��S��!Sw���	?����P0�"�U�ܫ7{ݡ�w�j	Ũ�
�9BPu
g~�����,�D�`��8F���n�'�Pk�u�@�g=S�֋���yB��Zh=�E��y��c!��,`i!�s#E�tޯ�Ð�^#�{"�J�ɽ�T�!��NC����a��4hX٥�R�|c�u�=t÷-�`��w�-����JL����)@���L+��(W���Z\X�3�K��VJT��8-��/���|�(�s�
y?���\
ya����d�� }��I{iʩ�� �0���r1˩��~�c���\oI ʟ
�E�q���3��~>�JW�m�S|�[baެ�oᯨ��p� 0\E����2�(�}�n�$xh,C	2��7���.�Q�|
����i�CI>��Q�_����L	�Ab	�)J̵xb���y��O�W^J�~?�7y�j*�j_M������[�|@/�H�)�,�~rW�?��Pz�-�56�2�H~^mx��[�08�HǢv�뭍��U�����uz�L�Y�8�f&���t�	����;�'��3��%b�X��#B��a���d��_�`�d���l)�D,?��Nli���0�z�s^5��Kx�(��N����� ��Q^�ZԠވ�l��L���?���^��:��`�gy�¤��3]x=v|Qa��H�~�Q*>g�'�!�3��J�����6���\���1��BsA�������0�ח��[>���x	k=��k�>�L�tC"
`*w� �j�tn�Zi�#;zĮC��+��X���k��O�z���V�	�I�L��ꯀd�2�1i�m�v.y/���� U�I��(�XӺ�@���R�]�����53�����Lق�aIV��3	��]+�e��=r���өb>����_u.:~_�Ѧkqc��p��[���C^��¡aῴ늬ٚE^�D����1��fde��g��2 �B�x_���06o�����Y��b��p~��]]~|}�H̋�1���[	������u�H$�c���q�p��l��G�[l��&�Q�CoE�����L?8\��al�������)v,�w��Fz�%Y|�h�4`kV퐛�;��4o�a�ŏ��2�$9�,�4��1�V[8�����7��B\Nӆ"׉���/��'��M��d`�Q�q�VΜY"�����|������F[�S5�xU�%���������8r�� ��'o�89��V��q1��e��t���6�N�B�)��-���Ƙ�'P�3�oq
u����=�,io��K�I�D����4�9T2X��(��|�c����=m��bU��k
��f���}^��,MGP7�x��3��v/Y޾�G�k˜z7�[Ƥc?���4�z�.�
WF������4$�_�����#�r0���dK}B��g⽥� �#�m+�xWU�ZY��;��gQȯo+�����
'\��X���Db����K6�c�75��}���ħh/M��ܾ��nx�@���Z9�LjV2L���kԆ��w�"3(7{G3ATMmu��N��wFKYGaR�o��b�^]k��8hcfG�O�y���/F��j�ox�N!c8RJ$�H�;� D��!��ѐ��#��4��q#�Q0S�>�*�,yX���E����N������(�;6�!���v�@�"	�`5���}e�5������~�km���m2�+��q��4ʎ��[�2=�{��O��ԅ�B=���e�";�7d��3X���������0��K���	�~���w+*Vg�P��1(��$��p��!#>��[{�����YHt))ihcª"�^��դ��XDb�jv�|p�*H�����x���H_��V
]7��Kk7o!/,��P��=YwEf9))
�#+����4;�?͵[�n��h!#�f��_1�s���� ��-�|��=���y���sG��Ҩ|�b崄�_ؽj
~�3g.ΊG^�s�y��zn婮5┮�w�D\2�ٖ��a{��8�I j�w�u�Dk#q<�4cҕ���P�B�HY3��ɟ�xg&���vm+T�kl#۹;���x�i�� �a�p~ڋ�ϸY�ְ�����F����_bo$��X���ય]�0����R���)	�Ʃ!��0Ia���(����9.��`Ǉ>U~��%��a�'�wo���O���ԋ�.��vC+0�/J�={��g�$
-�Zdg!/�l�z��y���ڙ2�Wl��_�(�zw�~o�A��>5�f��R����ȷ���=��?�M�,(���1ӏ�c���p�'|�흨�ݏ����fü���ws�JkIPJM�CD�_�j\�-n�;����T�iqŵCF)Ur&����;�m�mp ؤ��ZϹ���Y}�Ugk�[?�5�M�b}������8�|�>RC���%������өۢ�_���ޔ�Y����}�l�N\H!�><:B7��Q�s��yZ�Xez���	o��,W�5�X�<�uvM0�yЯ]d522\s�|�Z?�A���C+{�,;0A�^��ʫ�'t��Ƥ9�2{㖰�����>7|"�F*�nѐ)��9v�
ʺ[�5MU�������{��@�;�����|0y:��ʞ���s5�ZU�`�}r�Z
d����!�ʾ�^���>5#;c���)�gM���Q��i�cm �AVcGff�ʒ�[�o@�,�}A���!_�*Ҷ �9��`�ܣ�A$;m� �.r#޶�HWW��P2�Rr�S��Bצ܅��KM�#��6=c�Boӥa��g���H1��茁Ĥ�(%���r�|�����f���iɊ�������+t�'�7ʷG�Dd�}�S20Ȳj�Ed1�+IQ4=)c�k�P��@4���Y�6}�L�o�/����_v�/$����G��z���>��Řm�t23f���\���d'��e��5��y�
�Įq�	�e
N�Y=�������@̈Hv���4X� �(��?�|f~o���o��^�>�;R�w��a����un^q��&hQ��	F.�|tP��!��[4�Moce+�+9HJ�EsI�N�M�,H瘶_�2a
�'jn
k�T���N��@�g5x0��E��/'4�����[R����{��QKG{6�C�����>IjKT���k���z�����mpze�qx��\��޼b����(��
f(�m�;��&_��� (�'o9$=`Cf�Tv|fT(��2��Mg"����w��%�6 �;��p#l)u�J(����#?�ы�h}�}���|�;�1e��:��L�M�Щ.<7�e�C���s��>��}����Qz+c����@a�Lc5J����Bzs���Y��o��K]M��]����i��95�Zӝ=H��}�i`���:P��&��p�ڟ�ƾb;�%L��o���(�`Z5���D^�g�pkѬ�eh��H8�*{߯s�tf�D��^�=qbo|:�f��^�y�:e������n����q�zSp���4>��?�)YN&%��B9��Y��%�}M��t��b�j�cl"�&m|�^��� D=(DN�w}������3���Փ���}L�8��8$[7z�KÃ0(4�#�0q��p���a���<z%y�C������h�!LM�`m�J�Ѳ�(! �G�'9���Z`�-/�7���S���KP���lbF���]$�nd�r?�N�V/uc��@�3��"|I�ߟ�&Z�+Y8���\Dw�ֻ�y�WgN����b\h�[!�9侤�GM�
�|]��T��{x���`F�[��!��y�n.<��;n@a�=�¡��6�F�G��T�da��'���jL����L�&Ѱ���5�l�Dy��ȡ}����-nD�<��źl���^K	 0��-��� j����q���eS�\�z�Q@���iT{J��?m$��Ql�ϱ�h�� 7]'�6n8<w��P�~��ލ)���{�	�6I�jK Ԃt�c@��6�w��W	Uz��!Uŵ�C3�V�D[ziN�.%�,�lP��������IhI5~V�ͨ�2kCX�S��sY IJe�����%q`k!{Od�Zٿ��0p"���S��D \#�?�K(������qp
�������{i�{r?�o]������C�F�G{*�bʈ�� {����U]�I�)��}��G��3�*�,)����z���ʖs�|�&�E�m��-Cݣ�ayM�[zfZ�6¤Mb�}BG��f1M���Q��e��L9j����wp�*�=�;�<nHU�'��e
tc	�0{�t�~<ɞ��?V�75r�p`-�9!Z,5,�Y|F' ?ۄ�n�>�_���|r��B�#���Ԙ�*@�:�����w7ꀪl��M����y�ۊ�:e�^�].���C�ڊg��|�/����n-��jԯ(�LE� T4]�j!�
�c���� �㐡Gf/~N���F����N�s�3��P�Y���@\l9`��聒oGF���*2�)b))�B9�L2�ya��`�k����2�N_��g[b�AE7i3ا���\����\�e
��J�R.�?���E-��O!�(@>�Dy�>� �%�3����p�Ck��L_x����o&ެE�a�k��>���=9ڕ��6��kO�͘3�rV�7�����ۆ�w��>j�v�h���;�@xa��9��.�>zs?������r��Dֺf��E��D���\P �CDH��3
Q?��*M���Y��s����y��r���LC�ʖ�
��.�I�܉1�\�o~���X1�}�]s��[Q������xSK����A�+@�M
x�`�7&kP���`�T���B-�1���m��]�ͳ�p�U���H�r0\L��^�_�ջe� �چ ���1�?�"�?���D}th��<�K���T�;��@�N�A�o��*ɲ�I:�� Յ��ny� @Xs�Jg��3�� (r�k�T�XAyr��+�𰒆%:��M��	���̴s����6�	ub%K~ó\tsu �y��	v���ӧ9C�w���Ĳ���vL��)?���Z*N��� �sң]d��v4�T�v�8O�$$Ʋ{B���`G�]	e&��}���CU�KW~@y�>&���j>�1b|чUu+��ڪ����UT��\��*	t+2xz!���n��.	|���R��a��賠��#R�?��_e�rw��?,�2�v�c�En����U8�����Q�N��;l��oUrC&������Rd�R���<�����/E���S�9�˴�����oi�{?}� ��ĭ�D�+��Bj�v���J{3������ppv8��|�N��%,ɏ���2 Z��f�*�վE�|����r�WR1�d����?�Ky�E&�����xű?�t���\��RN=��x�#���:O|��1|��3���/G�����W�+k2�e���C���Ð1J���?7a&�qEn�nh���_P�#��?�j����!�	��$@ �]B�h�r�D[��!��6�����BA�/��1�OkD�������/^�c�jYԁ��/����(�����B$���Q'^n�@�͡��Zr�#� 1N�[_�k]`[h�E��΂�E�Q�ô�m��Żð�lc��~��)��KE� �-�gGȲc5컓�����{��p�7��3J��`s���k���m�Wl�>�Z�*���1	�=�U�t|�w����bP`'��a���^���'��i!׿�*7��tVr!lP�[r�Nd��t�����à�	�I�L�3�M�H_�%�s�[��u�.� ����]lR9�ߒ�C�H��n�˥y���R�1h&��r��[H��Jֆ,fC���X�c�eOl�EP��'�{Jzo�����:�ey]���.��v��`N��fe��=���#��+��Hæ�HgGͺOj�����<�w�� i��/G�.2&�`���G��`HC�6YUܬQs� �m��H߻s�-.���D���7ryf*g������)��8Q��j&�G����i ��<UlM6�n���8?C?YD���K�¨��[��+�B�LE���;O�iP\Q���_ ����C]֓浞��B���#�ښg�׌�=��*(���^����ݲ�� \�mHL6�4�+�G"?�׉t��P�dLt��ѥzH����6Ԍ����3W*�3��/���ҺA�$�;����J�Չ� ;G�x_�����#EXw�K��r�x�9��S��:�t�����9�w�6;��f��t<j݆I�Hŉs'��u�/B�-���	u^�X�-�+9�u�%B�Į����k>�!2R�����!�Ή�d-���Z�*��:��+���X���к�i�������1���>cƊ�7b&�=VIM}pd�4pd�?�4��
�������yH�%���jM�p���%�0z�G,g0�FH��eo�����m���
�����ʕ${�!,�R*� W�6�`�Ap|��Y��<��{���8�
����&��K����.\U��
�p�N�U�V��n٦�� �_��#��='x^���t/t2��C�y.aS�ż�L������&w=F�%�W@D�@Z6��5c��> J�\Y�hIE�Оhr��/���!*5߄�N^w�彉q9�"P_� ��;6�|Rg����a#�� �ډ��� 7$�Ґ�ɀ��p����䗴����a���;��SzϾ�l���߬����m��mJ8P�oO ��9�4
����{\x.$�~�bw�9�n�LK���ȌHW�Cy3����J,2��0��Ǥ�f��
�U�e;yBR_����|"4�B̏��N_��t'��,U���3,�?���U�As��Q�u����B��E�0M��g���	g>Db�+����ޫi�g�Hו~�j�G���
�q&Tb>Qi���(v��}.��/�v'5m��#~{���	F7\��y�fb��F���\�<��E᠘'_�
���ު��S���wjĈ�z�A��B���0�x����5�<��М@K��h��4��g��V[����k�º%��s�<�;�<j�m��ST���2���,mQ|���]���j$��a��V��i����ڮ�Rm}�@_�R)�pzgم�-��|��P^�?h���s�� �P�w�XѼ���ג���i:���pn8�����ķ֖w��׏�"Nt�rz\z� Չ>�m]`ʾS3$�T�;�tg�����,^����OEe�� ��p�"�%o����h�nV''% �U|\��~����x���&q(����/ g�F	����*���Đ�*����WK��{�>���,<��,M�Z����{�����Q���r�{������圬��V��֩��Y.8&�e�>_믡� ��G@����F�謨���E��z������w�6ts���q���l�R[$��EεEȶ�y��o�fB7���@(R��V�(B, �������u�B��i� h����?妫�U�A�;�M=�t�uXp�2�����d�<%��}����$��<N�Ae�J�2#������zh�����\���n텢���
3� �q=���4__ŉ�
%�$�������A��`�²�G-���:��I!��E��X@�E):�Ub��s]�RIl ���:��*�Z��V1P�$"oU]�Q�os���Q�$��π�q����EV�&T�T�2�����^A���5�OO.��kQ	�Jw�GЏ8!EU��M`�58H����JI_�F�V@ި�סA�a��`�75)h:Vn_�u���Cjy���hB#�a�\����V�m��p��3��I#2^e��_��+�D'
0'5<3D����*��;��C����U� ߤ$G�0��[ ��(.)&S��B3V���u���3���=��K�p(EZ��A�R�����v�s�V��$�,*��n;�rܞdB�j����X<4�?����]8���i.�r_N���o������n�}�����ي0{��ZCunlJ�|%M��j*	T�����Fb���G�l�A'�H���-g�u�t? �i-:Z���0T;��d���t�?KS�t�J�~����v�q�3�(:V��ޣx���^�| !�+�9�.�K`��0����7���aN͆J]&�NQN��A�:`�<!��H���)h�5oLp����������r3�/we��wk��sJ�YG��5�/�t8<�k�������p�pM��w�P&<���\;b�'8�e���Κ}�����]�
��Q�.l�nٝ��uo?zn�+���U����o ��h&�wp��S�G�#�c ��R�fV�8wg�-��?� �W�;4���]!��7�a/��F(D�ģ�Y��4�Yް�e���
�ɯ ��3Gw�z���  h�3⪘qs�%n����]w0���1b�>����5S�~ �r�7�N�����ɔ_�PЗP���,�������`.��Q���HY@~ ��|���{\�i)J,*����{_{�]_哔S�Ī�Y��2=����mPD�x+�Nq$lhw��rĐ�׵���^:݆��{�T<Ȱ��x�4��5��6��q 1��1�ʿ��p��6�E��r	�\+��}�R��mn�9�ULo�KIۊe�p��+GH�4j��?3��1��0TO��F�S⥙> 1�˻�g@��V8�� ��f�pI
>t�].Dm��|�ŉDW��	afS�R�>is��)W��?x>�����J�i��hy[��o�ݱ�/ݻ����� ����nu"����JS��/z�E��Xm:�'��DpN��&*֭��}�{�����e5/��?��P��_�q��#�C'�`~B�}��`�O$�\�O�l;y�Az�=�ő�`꓏�'������ײ�]u��՚I�|�2:{1�����#!�}Ck�H�^f�n��@�kH�{��'X>��~�W),#���tAU�l�ĉ~[1V�7mU���"O��?P}؃�
�6���Y1_���h�=��j�()��7�ͱ��:5Mگ!<#�:�l��_�[ƞfTʚm�%\-��; `&�~�� 
mΝտ�2���<�|�'�Ev��x�Y<���99�Jlw��H��Ph	`�,h@5�*a�R�YN�")����f�َ!׻���}��T��o�`���>���*O�}�i�8�y�a�Ӗ�p9u�E�Wٰ]��JV�Y��ctdUdtG�E����j�3Vs�߳H����8iSB��N��n)X��F�0{��P���Uerj�&Z�s�(��F�M�|E�
�h�Kn��}�G�=����@�uz�_�����y��3[�<=]��fo7�h����8�g�(��?�H�!�}`v� f�a�/{�X�q"��#��u�s����<�eҐ��a�}߸| kt�{��}K��'�&/�t�z��*H���(��Z�R�q�v�R��@�k�/Iw�u�(S�($��k���
��~��j8���\��lN��M	���������ޞ��s	?D��O����4���Ϭ2	W;�)�s�^SqP8�4Ϥ�32*��Q&}�g܍�8G��F�I<?��q���>�U�Xf#��m|e�)����وCIϙ���4�Ǩ���6�B4{BA	r�:XuQ�`Tkf��~fr�b\y�0�/b��܎�Wi��n�t(ٹ�j]�L}�,:���<�1�i�Hp��='I�g���`.��/wHe9~.M�Kq(^���r*w���1��q���S����נ~@n����E�#�1���d���:y�`Pgl�'����Kߋ=���2���I��Dn����[w>#���J�f� v���m�é^y�6����9b����GDŀ�|I}s��.[%7 ���ڄď�b��ԩc���$��fr�Dq9��δk��\z� O�1�E|�9=�1`��:��U��^޼+Aa��ǖt!�˟��l���D��H�@��Z1}�,��M�6k�9�]�$M6�]؃΁#>_d�Mϱ'��l/}��߷�,u(��L�kP�.�@�г�.c�G�v������}�Ý^����� ��\E�����frUn��ta�+��G����',0�"�YXu}��%����J�{����˫�� ?��|�MnJz�[f���"لC�R$���t�Q*�@��I��B�8��R���u=�M�e��W�!8�wT��4>d�pp]S��(��G+���]��c�4�(�W�F����	���BI6������75櫨3ˤ�b��|(����	����7�i\p���o�wْԾ�gO��&�}#�,�~j�'�x��(���#��(]��S!G,m\�bn ˚5!T�' �MiPԺ�\�.*��꾯s@$�.
��.��v&y��-��?��H�LE�Zx�7?ag�[�}�xe̲�V�q�]����Sq���^�q�����?�h��912 ��~�+JY�8��zam������LY��pR��D��&<��n^����3�	>c�t��'�_���b:�-���	�$��ߋ�J�<8�M9Vvn���^�����+8��,RCLH�,Z���	e��ׅ�=#��=�=�&I��ܵ> = k��n�ݕ
|Q80
+c�D�:UL A��{:��>-"R�<Z������bb/9�%�ԺB��i��#y��x�ׯ�K��V����i=�"��=�A�Pq*��L\��~����,`�f�7�j�?0>s�Ң��{��М�rz.v���D�FV?�T�Z��C$P(����G	��LߟVS5�Y(�Y\����7P��[�(8��~[Ӳ��y]��K B5;�G}��1�2jN!]h7�cww&Y1q�V(�_�9�������)0Z)c�C~������Mk��*Wǡ�P���ӕw�'�ufa���X _3��M��|KU�u�����{v0�sq�v�W���o��������>'��x����̅��X�	�_�L�k������8��1��H20��숣"H]��jwdT�����T��8�H�þ��g�Y\�2������Q+m
n�/���*�}.e��2�֒%��3�/���芾�f�>�7�	�5��U\�I�j��C&���Vz�*|��d�7������̆����͡��Al�jiWE�^*�n���!��K'1�R�%�B`S�%�i�V���y؆�[�OG*tq����n�R�@�x��(�u���'�v��T�}ex�_�2�eʋ+UA�U�����M�f���5�m� JF�8&�&q[Pw���/\8ӝT�(���R�)��5����ل����.���S5o��3�ps�ԙ�>�D���;�Kp쮓&��Z���C�A��j��{uT��F�!SO�䶍@�̳tlT"��	=7��
��,�wd[L��n�a����q����'�ʲ`�n�#ۅ�<t�E#UE6qMY�.X�<EK*K�tN�f��M�R�l�?h��yk��kx��	z��d8qǏ5�Z�(47�]�o�D���] ������25���X`�J��v���Q�*�& �oZ$��ǧ�!�_�����Gf��w�/;�T�#J &�K��@��dwkw<�<��b3͕y�s�b��Ա���da��=y���@�\�!�3g⒟�#v�?^zjQ���8��#� ���ݺ�����}a��2�U���zv�3(�����}G�.�sV����xf�l�q=���I��=�&�4ߐAĞ�J�t/�h���DF`���w�����v��L�$�>�i�B�,�sL;�=gg�Z�e�k��W�Z/�����O��i���rwf�̪�uߣr.B&>��kH�Yٖ����/X�%�����IJ��	D�64�\Wl�U���UY�a���{5EŲ��9���>"�9G�	��U�z����`�bQ�ơ�Λ�����u�6��Y&8�%��U��"�#*���-#���;EE�F�8�h��jƗ3L\����"���ׅb?��IY��b���lݩ�u�^|�_/��4ĵ�C���!�E8x�t�D0�v�]�OG������u��F��Y���J8����ry���&>Xɫ�E��P�H�E/��:�
����H3?�d
�����z&����p��%���y���j�Ev�Z�P]�X�#~̘I:��S�B�&�d�f=�q�ܷ`~�+�r�Qj�>>RR��n��=����t����z�B�{1�ê-?�5��1ADK�xc�Zj�u�F=#[��|{kLh�|��^��+'KB3�m�e���h#M�WN�-�&I�OTj�� <J��wpA}m�t�E8Z>�U�/�(9μ�(tR�7���,p߻��h2*�s�y�^�5 �dNP�^12���J�n��F���ن�.-�Z�\H(������dL)�䝿�d�V�Jl0���-Ӄn�s��F�m�s֑���p�I[�-^Pc��}�<h���?u��ʖ�y ׷+#�5�r�$��F�_�@(�-ڧ�R�ڭp� y���
�w���"-;E����35qU������N~O_���6���*�����{."��������3��;'�u�D�}�p�k/��-�v=W�v�B�R���?I���F��.?Y�"��Wб-R�� r�	�l��\H�]	Y����#X}�Jfw'��i�[�|]���A����T:A��Q�� ��,�,����&Y�4*�FL������&�=����t&�t��� ����Ms��G�/%�㸾Q/��|�9Ht5��j��N�"�+s���%�B��FA�8�J����BJZ�"�d&��yp�e��+�6���]b�ǟs��@�D|䢃���]p8����*^0��u�m*��׹R\>�6<2ֆ3]ü�:�f����Ì��9WN-���^ڢ�LD��\ƽ��s�v�����?!"��u�,�)'�'���[���G)*�`{�X��_����û���E'Ջ�F�/(=h�2]#=�Wt��gr�:%�*HY�栧}L���ؽD=p�EN�s���oAo�s��1$��1���}�e�}��9ﱀ��q깹R%v�̴1�,Fϴ���	�B�F��6��I�w��І1���->Z����!{#0~Q����q29�B��h�H�[����k��g�Ԅ��m:�U�(7���%�|������4H�ᘍ��'`�#�4h���?au�a���8������^���㊡Xd�Nhi���s-�ڇ�c�n�#fT0� +�q���'��,(d*��}���zA�B8;�u�T�6���P�dA�$,\׿Q��>49g}�GmJ9+�+�^ze�D^��ʢܬA:��.N��߮��?�j�C����G�«黜�Ǻ�xGg�����Y�����HK�쟞���kDF���_��A.�Eȿ�=����W{�,:%>�}t���ρ���ƛ4��ږ�FF
�W�UU��FK��o�G/�ظ-� (1�R��^`�0��E�YY<�߸��(l�yӿY���G�#}�@��~�u¤m�PV)�=��[b�&��*�c��\���!���w��߻�����'5�*�'=�<����ܸ�3$ݡ�����`��"�AB�i[��D� ���^�e#-闉#�'��Sj�f�ye*U\u�ea��1E84*6�6�p�XB�1��8{t�l��½���R��Y& � �}s�]�r��p�lq�
�	�C�gl�V{�&z�����|��o��i�R
� :�@,��y ���ie�77��8`3�q�q?z��Vn�z",`I_��ة]���e�7f�o|�DNSj�q�GJ~/��4��Xq�i'�]%(��\'�l�h#z��{(}Ȧ�#�	���Q�2u�a���5�UJC-Kal�g>��*b,,d�F<;ZR��Ih9�<�h��ی$����l�E�a/�nGǿ����a��J�!��a���J!�~+�-��XTw��ɮ�E�~R�պK��$1բm8�eUVek��&���WACy���*��/�[	�r�����F(�Xl�r��&/�p9"���i��E����B���p)�>|~�蟋o���D,R[�CP�k����㞧_'��v�{�&&�9��3���o39����g�/	m#��H&6����X�H��A P2�B�dm�=�Ol+�ϲ��F�dW���B��;��
�+'s�u(0l�4�@<���% �N�^_�- ˴�?�;�;B�'B a���}��t#F,h�9��\��Za���-�Þ~y:n�<�=A�e�L�@�~J�P/^�J��<H#��xOl8+��  �s�Y3O��1�B���|T��{AV� ��{�x"9v��A -"oG�y�Y�31�դD�	,�ʵ�i�V�YK�����H���`�%[J%�*��h�a%@P���|����<����#E��u;�5��EkX[*��9�UG�)��iI�>�ٌ�z4�w�W�-��P	�npYF����~��6C">>0i�ߙ)M�\���ȾT���~m�Vݵ2�#��9tJ�i0�-bI���]�*�~gY� ��i@h�����ZKN_0>��9��X$W��������1��:���<S�J(b
�bM���еKTcB��A�O"+��q��B�[�nQ��\�A�25���KH>a�Be�wƠ��~{�0�4i�W��3�{�Mv����렖}
V�,�?�sڔ�o.ݶ�����!J��EϨ�;D��J�H\��������8Ԏ���W��b+'ﳩ�i>韤Ƿ>��R�.����â6�j吰m&2�җ��sW��|�W�/I�4k:v2рV�۟-B=��{3�c]7��۳���P��K�����D�گ&+��^�na�f��|"Q;� ���)Ԡ�D9H�|c��|�&d�H��"��Q�wY{��p��~[ʕ����tH0�t"մ�������3~a#�b�#�L��2����E��q'�5�o�o�V�]�Q0ZV,�t#�`Q��Rƽ�h�d��o�p�]A>�����"9�LMQ&d�#�6�E����5�.�E�w�d��������!=�y�t`��/Yz�䃟���9�j�A$���(���A�G�`��������ˋ[�qb���j�2������X*#��e6������o�\Ɠ��?�(��49�'�t�N��~?^Ň�u�h�@_��I�}%ԅFrE�f���b��J�[��G�"S}^hxՓ^�Cj���g�;�c����w��_��_�jY~о��z��%����gԡ��,۲���n9�b����;��Q� ����@u��]���ӽ8?Q����N�h�m�g�g�B@+�@rU��m�u�"��j��s���Б��M�8��p��l"����l����y:������t#�Z�A^	w�m�ᑜ�䱻Ʊ��%\�j��͑�z,)�`4M�l�,}�4ˎ�wuOZ�ɠ�a����9��Mvܦ�C�	r���}a9[P
5�;J����!m.B��C0[�]N�o���i�`%���Iկ+��dׄ���HMa�ε�)'T:<�H��%5$N�_ �\�d�|[e^L6��?�aK*�L��mm@R�`�56��ͩsed٢INd�,ˎ�gzFp�n��O��Z�н^ɿnb�h��[׵�*��3n�L���~?�{�Z2��>l��>�}�+W)���$��Ѹ �G^Y�G~SsX��H�l�5�l���E��*�;,	l %�Ǐ(Y�*q��P[�4�������ʻVDu1�pKFZ��aʖ�i�C�Տ3��� ��� G�����Z�c��v�Z�Y�A��r�ċ���8β�K�n�$Z���mM��{FT�qx]����QՌ3,��0�o/8��:���WyU��m�/��	3�(�����ˠ~QR_*]�+�Am������W>V�bZ �v�.i�Ey�?�+A�ThC6����*ٛ#}�Y�`��|�V
)�IG����?�i!�!*���] T�ˀ�M�0�4�̔3e�>���t۰�)�l��8��u�I���l�t�^t1*	 u����^���|�b�K��X���K�2��ޱ,�o!���Q�<*\"L>�S�@�8��vņ�˒ϋ�G��`v@3�瀸�uW �~p����$������#��(�b�i�ENK��b�I��`�G�ޚ�p�D��.��<��b3���{`E֦Д�#E�D)>��v���P��U ���`��F�$�Ri�*�I��x��+�Nu%@hizh�,���&����G;x ��P��ғ��݅]>�-���P5��,�K�g����{Tk�e@��g^���x�<��rο}�"�N�?p�
���'����&�����R^[`4��I�n-��K�st�J���ʝ�YĨ�ЧvS���xeE_@�Nc�Z߭E]��@y8���Π�rB�;����ǿ��!p�-ms6���f��D���Eįw�'~|�#wl�w���	a?��*�.;d������$�9�X|LZr���.8���Yv�|<mjAԃ*w��G����[���N��6X��Q�l]�K>�9�XN=��)_���.0���اk�T�2��˴�6=����즓@w��;��Ў��8C���r��nQ�"j^�^�Б��Ni��8mȡt���Ngph����B�r���&�?����HW�?}+��#j#^� �������l-�_®��h�m�Cǣ�U����P�;�����+j2��_��ݒ����4��m����@P�"i{�<g���%�C/�#�E[öA���ȶ)r�>HZ��AOt�fݴ)�&@[!����q�"H}�T4 �=��d�M]�M}kE�6���y��i>ӓ���2+|8A���� �Dڲ�4���Uu�\E��Pf�`��"qS׹�lz|�� 5󎂾�����Ȇ�(-�ڻf0����HYB�[X�c-��t���C�P~ss]ή>� ҡ��/'f��|�)Mۘ�T�����Nٞuv�-ώgIL��PG-���w��#�{Q6�"lࠇ����?vL�gf��(�����Xs��9)�l���� _.����ՒN���۫
l�ؒ��g�ܝ�.ՐtYG�"ˣa~��{��*߻��^p.��-ۛ�M�[J��4����b^"������n�*�~*ґR��K�+��:,�bo���M�;7��CY5g�.�Te�R�o&Q�W�a�f'�������S�[^qY�LqG(��k@}C��/�i�X���F�q$U4��$���Ɛ"Hj#G�G��\����g�R'����6T�^cjW����|�v�rM;�M@�P !a�ɉN�l���k��IJBz0/2���Ӛ�}�iJ��w�9&	��٨S�ߍ���O�d�j��� �?��X�W�'�F��O��&��*>α�br��$$��wY^X5�AD�3���Yj�OA�}]�����d�fҀ�g��EܜO�e��p�׭0�H��Ŏ����~� yv(���#H��{g�6W�%�e"o���b.IX��Pw�罚Iاܤ�p��L��E��`%yw�����P���"0Si:�@T|	B8j]�4z����p��s7�B?��{l�m�;�$���5֩p+V�%��.h;�;��"��욋�*pKEu��,�YzD��;s������GQ�� �)	s��=3'�w�3���R�����v�!ۂ�/�{e�6����C�&�Q�ķɬ@%;b&��N���
3����_�'�s��m]A��
HOGG+!�=��l����_���МH⮖7x�r۱��.Y�Lf���0��O(�	Ӎ?I�+@�sG1�����x��{��Go���Du݃�Д�Z�1�y�'7g!�II~�P���k"��:����p�i��0����5CU����M;���QPP�mo��C��������ʹ³Z�u��L�H+�-����9ղo�&��2�j�z\�r�\Bh��=q�T�Sό^�r���TZivn�[ *�0ph�1�W�]��~R�K�Mg/�����{W	���I�>ċ
�֥�:>�>�TP<uJ�F�ȍ�qs�����;N�1��F����f]!�)�[1���6J�w1jhhVj���E]�;���#��w�qb-�.���\�`����ui�k3	��j�oO���]��",���;��XB�Z�(����!����k΅1��:�<��2\����~�;Ĝ�~�@>���+S�G-q&������l@�~�׈��Ex�r���� |'�{���=nX7�^�(��h�"2oW�C!��o��t�k��[�[Ѵ�f#� ����4(U��&�6��H<�:���e�3-�>?����N����UA������}9������J�Ƭ�>����45L��-sj����Nj�ѹ��.`'�&��_�X���Ca%B鮴T���?�$�/�+���H�����Nی��"�kF^0��u.�����F�_�*�S�]������T�W�Yd�)�u�҈�s}��^G�Kq�)�OES���^q8B=�wu��i\�;r��y��k���_���8�����9�t�Do4!Jڧx�����=�;x�J�Ʌ�5������T�C!�DZ��c��Z� �����\9�K�mC��4�A�0t���."���ꤑ�����%����ĥP����/��躅Z9_�^k�H<�H����L#��GF�4K8D���`1�"d�]L.g_\�r�|e�o1/ʘ�]n��@/T=�˰��ٮ#������:�;(ծxH���WdO��e?A�ݝElݷ��O(����|&4�s��\>��W�V��HIJ�+���jl�#^Μ�<Z��,9.y�mgƇJ�U�N?c)`/(V���� �N
G�+�h&A|&�a�?؊����}�"�W鷰B��#����'�RR�bJK���냿pv��$�ɱ�U?ۄbyv_(ȗ��+o(<��	�Ni�#xy_��D.�Z�z:P�W� 0�C�F/�����ٺ��g��V+�ԊY��DCA�T4]L��E���
���_�-��mo����d�x��t���m��sw�k�����!�g�f�����vr+�@��	�:��S����3X�����.RW�	���id �]��ӤX��~�U�M�x�)�"�YjFٰ���O���W��T�,��>+���eW8}˳�Ϥ��m�WN5�v��b���n�[�?�,����QR,�Y�Q�|�n�U8�A�T���韶����LX2�ԕ���nF�o,}���Z�/��4y�꬟"�/B6�� ?]�e^�Bl�(dE���ZK�8G�d����@���=J����K��NC�3�`�B��>�;�!�[�+jЩ2�k�kB�y�����)�5��\��e���Un��h��aT*QPIU�1IBW�:;�@�	"�14|*����}��%��!C���m%c}ӻ������j5w%�x:7g�´��F�B�D鴻�VMI�qfx�b{�b���²0��6J�����HS k��z�,����V6q�#!�CNV(�r �r�=6�e�e��f�2��B�f�(�C�A,�����N8Y���L�Ԡ"o7�_�:�}U
�k`���Om���>�.-
�W%����֛������S~!6�u�������u�����|�$��?2t `^K��w�a�����-6	��ft�!s$$�c�]L��4u	֐��W��d�u�6a�:K8�=R��g��(��AJ�U�~7��i`���?w���ۼ銪��6�.�#��Y��hF�۵	R�5�U��O��pی����~4�����%�[�~QU�QԺL;�au�r~�w�XǺA����b{�����UO�$�kL���>�P��*��5غ��C�v!�U���Gi�`�Q@�m��h���x�S�v�jqW�ԎFLp�������� �[�(�V�,עZ��ֽ�u��@�TW%kb���H}.9��� �2��|�(
;�|P*�	�P�6�]�{�������6�����p6jt��&�E��B�`��(F���P�2Cn�=<Q�G3I��8lg��n�,����e�;��9ȥZ
9��R.v7�#OT.�	7�lH����}Y~<�_�()V�������C����*y�UA1 �d���A1>zg�$	܁|�[�Xä��[��&��'6&χox(��̴�J #o�,��՛��21�}qk���Jp~�7.NoU�[B��ӷ�)Gs�*%��=T������2��4�Jm3T�۩/�g�l�B�]��V!�
G�62K�m�+�ω]��zK�����e��`Y�v/'?X\��P���p�Z���E�-�����;s,?kB�[�63%�����B��F�mCdLw@��zy����
A@!���YPw�y�\Hx���I�BG�c=���eh��������.��q��N a�U Q=eŖST������oB����[;رT�k߇9���3D`xѴ(4S�$&v��c.��g�����~Wp��ժ@͎���HГv(q}�*]$��v���+ոht׺o��[x+#�AA"ϲ戉����<�I�DM)$���I�_�xNX\�yY.}��C�~�H�z-}��i,3��a"��_���+\��(O�]P�j���������$79P�r2�y�ߠTP�pJH�\�FO�O���;-�Ƶ���W&���*���e��`_R�&�1�#t���S~�7(X[����UO7dUC�~�Ň��q�l;��O.���)b����뫍�\�R
3�B��uٙh��;ª)rvP.ϔE�8ϩ�!�J����g�ǰ�g$�L	��0;?���*��#_ ?�/��LZ��_��\ߋh�̺Օ����
��Y�5�px�8�䳕�!N�i����s�-�(���ȿC�/XT���CF�M8oS$��'��L2d��EA5���D����r���2��mъEKQ*Xh�Vb�CI��E�y�����.;5���P�m�2c]kX+�3k?b�+�WU�(�P�_���#�ޮ�OV�Ŗ_�ǜ���B zÚt���P�hV��t����R��������R�������RDZ��jh��=�3��K���PgU�q?Qآ��s{��	����@E]��r�Z�����	� �)�$b�*�f���Z��3�jC����qߡ<���=`�y�}�o�ʑ�����]k�޼��1Ӕ���9ʋT�ה�����)�����5���j�%��S&P����X��N_�-R�c���9�?
n���/�Q��A�{���T�M�+��V
��'�H�m{:-5[�"c5�r#E�Ʉ\l����?|V�c���愤�O˿d�_�jj[�𘨥�~�N8��)Y6v���ʓ���yU7��%��_�u�F����M��]=d9�;�ȫWT�� ��@�"����Z����~ߘ�U�D@Qn�k�6ޘ�� ��|�l��z�|���͓���?�p	*��!z�Aqg�C�5�T�N9����%�N���B��(b�������X=�QH��}9�����]|u��m���~��q����n��1����o�.�ˮ�',�'ٹ��v�UX� w��x�h��[z�΍�Ƈ��o����"|߳��U�D�&�f�;�}� 5����Mw�*::��>z��Y�IJ?$� ���c�t:�v��I�d$���t�a����ι)�RZ��z�[P��e��8�	�����;,	�>��^�U�N+�q�nZ��'˓���D����F�l�Gp�C
�a��©��B}Y�~7�	�����6����&A�J�b�O%;z��IA�u�_��(�F�:�"(�L��WM��(�1��DJ�٨"??��ҟ��;�=�&q�vq���v#�=��������ܛ�`�x��
Ę�on�x��=�*K������m�lK��6�̩Rfj�	�8���pb����C �g<�������Rl�f�x��9������;��������<c~��<Q��ĕ��YS�j��g�P�f_XB��"�>D]8�<�:WXy�?	+`;(�����?��S�t�gKE@2�u��7G�z*~�)}WL��!��Q�}���g=Y�v��Yk���Rs�c	���Z��J�6^2��������k��a��`S�.�4;Q�Lsd'���$�-�t�/�`���"H�v�u���UN���B�-P%�E
���w���S0죦�W5Vd��A+����m��L��i~V�ZC����y�f$co�KW�����O� ~�z*�]�J� �8�س8 �j�=6S{^3�W���z�=`z��~"x���D	@�W��p)��$�w��Yϴ��(���{
�;(4k(�%���L?B��4��?��[�S����8d(@���8l�=�-�y��+T��*��,L�y��ޡK�aW���E�l����𹣴Z�a><['K�����j���J�e]�]!�69��7�@mU��:8$퓬�k�Шp��|�������!S�|؊�׊'�8=�zp�O��"���gL��~D�{�5�����JK��y-B���&���l�����5�6m�c���vEޙ�lؑ�${���s��m��-~�j]���#kmBklh�Pxv�Q�dߙ�fn��$фI����w����e֬D~�1��Ћ8�ꔗ���-'L�nm�p �w�4�e��Y��Ŝ��;>��l�q��� �6ra���� #����J�lb&���_w�h#(��å�Q�Bߨl��i	`�n���r`�����Z���'>Z��F'N���@5Z�&���K�����F
�F�E����yN����j\:MnU�0&�������h?��%�����!���W®=���@��ϴ�ԲROF�K-n�*���<��h��5�+��ğ��w}�������i�����Ha@[)<���@;���1�����S�{,��B M�K3�q�M���(�����V[�˿���9�H�k)��}}��%�� ���c3nɭf��S�y3��_\̾Ѐ�����3��k��/X�������Ր�di{��Eh>��h��gK`��A��OLmMV�
���\��U�v����C��mf��V폀KA�v�B�Ʋ'Ϻ\X�zS�yV���K"M!'�ΫG��]���L��f�H��h{4Q^w��������|�)ޝ��ɮ�A��a�'F�N�1�VPQP漀�4Eh(-�3���Sn��h�t�˗vρN�����C0ױ�(���H���؊�̦a��$XѮ�?Bm<)7	�:�6v+1(��U˳E�k�I;34|�3P�}1�U��e�%��56��'y�:	f�zL�rc|v�#����s�/[?��т���M84Z�y�/ϙr��H�+ТT��\r�Gٹb�rhA]3*��c)����+�~	�G3�aR��Z�ԦY�����Po��i ��!r��/� h�\c�o��"�Ϯ*[,L>Q	�b�5��O	83�J�-������,�}�]j��}Ŕ&�*���ۃ�� ә�C2�Q\T�s���[����Q��AL#%M��Xg�^2m-@!���/^t�ȏ|OQ\�aN��lt�@��.'��G�C��K�l9�8H��lDn�<�\?�L�a��1af:����&:v�Jx�,K������A _T�"3m�f͘l÷���: �0Nd���,;>ĥ0�O�j������_���?�]�~׀�d����CJ�%���JϏ�ѨX�G����)����׀�A�1�'�$TcK9������������˯��G�G���wJ�W��e�z;����{b{���%tJ ��Y2�=^�Qwp)�9m����5��?۹���\&Ǭ�8Ƿ,�P��؄s��q�0�>��<84c+h����e�O۠J�(�43�'}�GA+�øK�S��5 �3�;b�������n8�R
��{�yfL�3Z7T[�X�q�ՕC_�J���Ԛ�`#ɗ~�rq%�/}�r��id|l���<G���/�U����,Ʈ ��(9 �k<���=?SK��T]�+ɓ��e�dU�-�����Ub4	C|��̈́�T��xk�)�IGe�!+Gߠ�<?_�(E̱3D��D+���@���isFq�E�`���IwAC�
u��!��a�܄����5gO�]C�7m�;����q���l��n��h%���Q,��[ Z�dB<�	L5�*�V/�!��8$d�D*��o��u�ߣ*&�l��e��m�~U���X#�d�٦VQ�8�U�?���$������=���[�}��~[�ՐZ�J�Qܛ��������EB&�@��ġ�Ң�\𳓿Ǘ@J� r��cs�"/���ٯ�uIJ�&�/�D���z�Q _�5�W��WٖT͓��v�d�+��A�q��7��.ky���O�I .��P�1$Y�ق�����@����RF��&;�y2��kZ�P�2����/�Cw�wgƿ�୷�a��vVplX�j�`=�}@�62��K����]�X��=(L�����L��J��@�YX�C�J^r�y�[�Ӄ�u��'a��T*��n�
��U��WE�PD��(��k�ŶH�ϊ��|�a6*�k,��i�;u�Z]��-~��C�'z��E��#� z�l��\�m�����t�P5����_����__�Ϳ�C$���7@�st#P��){�DmݗP�F��g��_l���l�|ɬ3����I�W��,�Q�h����0���#
%E;vw�T/��ѕ4rՏ�9HۧQ��0�4zt%��A旤�(-^�y��NxR�2���0\)�g U�sM�Tܣ&[�c'Fr�k&l�m�̏67�����кA���:���M�R�f�7��GZ�$�A�����8lRB��{�q+C���*�z)�{w�O�R+n�wc�q@^�6����_J2�� FQ6L~W��,ǌ�k���e8%��ّ B?i�"�|�iӌ`"԰�\0e��?��Ό	�e����\ԙ�V�4>���;�|*V��k���J�+jH����iYe�/�)���Y�3��x ��.���t�ƻ�ɞ�&o1��tR�5P)̖a��m��'bQ��Z��x��s<h�/�����}DVl�^n��v��fnv��u�� #_ٔ8��]:��+L���Q��-{��nw))����R�}�"��F�Ju�%�3�V	�4}Z�ѷ`)�pg�m��ų�ΐWm�D�k�\��N�b�5V�>����\�TF����u=h�m�K�!c�go�j}s�� B@�R�R¨�� k�k��k�er���z��wK��r������^OQ�b�4�3��e �Du󿲠�[41̃��%�Ey��5��D����Q�d�
����VU21���gަ���	E��ߚ��'ݬ���?��tBN�0m-�^F��X�`�uWLZ{��~k����l��N����w�f �e�k��o`P�^��W��N͔M�׺�峩��<�I܂2���cuўN�"6��������c 9�g��Kޱ �1�k��W�P�����s��q��:E��C.+5����o�^�$F&%}����8f��X_���D������;��ԕxCV�򕠈>`|&��Sت��z����L%��xDb�6{�
�WQC��r?n�(�"c%db���c�����3�1Lس/��G�̺�I�me�N��HJ�e��]��}��,����¿��wZ�~���t�Z�ʪ�>�;I�|�*�۽�����.��������s8J���*��E�<�:��Y���|�JÔr�.H�-G������/�m�L�\te�E����V�w�Q�+L����O/�8��������o~\�6��_nΠ/Z-V{)�hU��?��*-|�E9h� ���&�KNO���R�%���y�×��o0_��u����.=���ݒo��Q��ͩ�$ˌ����v�M  5!���qcu�k��/�rX\��*!ޮ�o��H��	�&��pS欚Pi>��Bd�m�T����U�g�$�����iZЎ�aF>�����k���y>`��KL�\tcD�>�g[�2�><+�!
�\���r����I���݀��d $��1!�i��;T9�$�Ef�o!n5���pb[:�}{$����ITA�	U.��|j�l����ИoT��vX�X�jV�B�a`�QR\���=����K�_UJP#@��Z��$!d�����!�O�f����l�����_���
L!�k�|�4���.����Aa� �`�Ǫp���T���P�S�"�Rt���z����n�����ə��-H��1��0s;f#%F ��p$�҄y�Ж�J�뼴��<(!�����A����������	i�u�(j�RY�n�"�8�h�Z�n�!g������l(�`�>^1cV�>���%z�+�w 3B	vݏO�ά�0*N�f�� ������)��x1���˻��&�u��q2�a�aP���IJ,��Y]3�=����'��;�<`.H�ҹ��ީ��AX܎aq  ں����n��������A��~zm�a�U%�ߓ*l��3�W�ڃ���. Ɉ���\v��!)	h���C���&E�2�?����m����o����ό�[�h^�� �g+W=���E*���|d?�-�-�V���C�6�J.��_��	�����g�pȨ��:j�[W�Ș��G��Ĥ�iy۳J��By*�Ⓧ� ��10P��A�� �^s�㔰��Ǵ��l�a ��ׂ�(ֽAE��*x�����+�)߾���N��W��S-+�D���	4¶�D�fS�t���P�F�T�ozih�|1�T��A����(��;~v*��#�'�=\�+�.��j�������'>9b�B�zMYq���c ]|ڣ���s�8��VQ����M�uğ:���4g�C��g�_�Fl����(��o
������`��=�rėG����`�����b�.�qHm�?�*Nu~G�&t�v�7˺2Er�&�Od�\���N�n�i��i���\�8mwz�(���x�ۅ��"_��'{����?���	���5�>.�-X�%ι.��r���6�Z��f���P0�WG�_5a8@K��<�LJ6sk^6:1�=2AyI} k %БIO��������G��E*Gl�rp@H�oA�kU�K�O�\�o���M>���kF�&m+ئf�|��J��t�4����Z�_s���I�kq��knL
L�h�!Z�V�H��kWƼ��V��5��Z�,^eZ�sVV�?;��o��e��Y�(75 �0\��2��Qz�\�>�
x����9��c��&=%Ѭ�-@8��i��f	>��R�r�I��y!�c4�X���>i��=��kH�2���TӫZ��[_�,
@fQ�ʉ-:��<��DQr��c��궂���R8�����U*5�<������ǻJ�2Mh�_k�$������~����o��iĢ�q��\"8�yiDU�S�; ��A��|�-�c|�����뿾(�C�5�c���"�
�c�I��|1yR�T6vy�XP:0+��_��+Z�DN�H�}bcA��T?�\b���1��7	�w};���S�C*Q���ޮO 8������IX��֤v9*�I(�]~�AZ���u��XWη�W�Z�����$�L[���9#b%���:���0� 3[�X�圐�;���I�F�}��B*���_��]a:�yU�&z$U��O��x�S�0����w۰W��óT�W��K�TRS��xcY�ʻ������O�q�[#$��z$')E�!���9�8^�B�o�!o�D������>�g�>��ʐ�}�dpto�Sr-���E���E������qv��j�B{h	�f��(�,����&�T�k��R���<���n���Q75���+�9F����"u���o:4i�7������IR��D�H�Y�__�H��6:�T�|����=�b���0����?�Բ�UI�#t�m@�z��G%��"?X��K]��dˬ1����tf��0b�"b��HD�}�g����� ;!�fP��[���XV��攢h8�y��ȟΞ���>j^
>��}O~xM䗹�
�Da�ݥ)�n�o��[��[���۷��	��x9��x��ꃿ�)j�9��Xӄ�W�9��`@���oWa9��,zҳԘ�@;w�mM�}���w �Hi�^/�)��������(��"�ƮPh�|�p�zx��ol'�d6��� X��It@v����)��a�A(�I[�_"��$�i^P�F�L����f�0��E��֬�`��:|.0k9�tc�X��tm�[�]GVd{�̨�X">���|iK�]�g��ߋ�otQ
�}�鬊�R\�jɴ���p����_ģ�����@�}v)�o�~��`�NV���"�/z(p�/����K��q�A ?�F�·vm�-����#�
��e�q%:�ݺ����ԯ�X$S���V\�_G�{ӊ�l.�;Tt��e�|j
UT�}���5�?�v���׭���������E���tq��dN��!��Y���k?��˱��"��	Y�׸��-�UP���+L��Y�0V�Ր1!���_G +a�YsA�Q�׼K�E�ۨ��WU(��=!"cr�@C'Q@��� ���AXV�5�6�:��U	��!��R�g,m����>�hf�=�14���=�T@��������|��y�t�}���z�Թפ�p�W�ٌ{�a�n���d����գ�CR�Zh �M`v�턉�X\(�d]�����>3Mn5���H��B>��L�?��Z�4ܳ�`B�G�/�e)�b�ل���x�����ԄN�aQ^���h��g1���_��~�L�Z�-��oK l��� ��AJf��YAH�c2oSWLFz?�ŧ��f�a����a���I��hB�pH$7|ؕ�w$��".�~�u���Re-�T� i��X%R����9J-ptA�C�5��
��]�UU��a��M�Ҍ��G0�gӣ�ZBC�t�Q׶�_<��$4�Q��R'%��򐦪B�8	�t���ڑ�C��Di2���k=H&�6�NT��'wC�S�n2m,%�� J����ڑ�_��m6n��.�����ܴ=w�����naڙ�w�t�*׬���{��¿�H�+M�����Sx�j�+����c��m�02!�
_y�qWA�������'���Nm=L�5�ɣS���Ѩ^؃���tB�����Y�IJ��4�vZj)���LJ�ǯ`^1mhYY��=���n;V��~���
�ңU�~�U�3��x�i6���&q��D0�Qޡ��Ѯu�d(�dXɜ�~���e�t���������MԦD��$'C��Q���t��U�-S�۔.���W��vK����(���Ϙ��G��R0o����.���H'���^�S֒O��9Q+�6�[\ �q(�Q���y�\�D��=V�VD��{�E\WJ��ԆE�ۃZ���Y���[c��]�};�:��[��npt[Z2jJ�T�~r�$P����M­A������Q�>	-�å�k��f�F�񁏑��GR��/�B�8��w��\sVɋ|��~��'o�ۻ=f� �ٕ��x�Bz��	6�~�zd�3n�tq�����f��D�}����@��)�z��>���܅y�=��J�l�S%��qg�ʜZ]��
I=����ِQ��������%�U��R��������#VȈQ(ۿ>ǻkwx�i�fV�Σ.�g�tB�Ѕ�.���0af��Mw����
�K]4�����:�?\���kȮ��*���D��;���+m�E�.�z3��$�"�~��b��G���;82�^M^��\(
�?r�P��e{8/���b�n�oO�XP��"c�"-����G���`�
��I@&�`��#[�f�����t��@bJ��8�#>c��(j�0���n�iP�t����� ��VQ�ym�k���D�.d�2l�EU�[+�a	-���s�r�4>$"i���_|Oٳ����9i~�"T
g9�*j~OӪ]A��;/ق`~��ە�����z%% �h�YWH�j�u����7#F���y\���hq�C>xM���Bz9�HO&,bb_!m�_���C%���JD��uy^{F�������-�..�����ң�R��\K������v���+D�l��N���Tq�3����?��+��:�{�*).I~}�o旯 ���`�?�o�*��|�=*����O�R/�2�G�&/���f�K"V�3P�or��`?��;�`�� �7a�!U�a ��L������6J�{޷�r�#p�Td�����4�U�u����`��o>��4A�U���7wV�78T��)�
|s������{s%����Υs��>������^�fX_�H[��_�e%k���m=A6��m#���3���}FbX�!��!�}�L+���H
?��)o,W�y�2b��-ؾ����k�#�#ʔ{��,c�1X����#%���#�3S�(wQ*ι�*9]i����d�`�G�`���D�g5Oo-�;��~h���~�wՓ,�U7c"�����W���@�RλV0����x�V��1,ny�7����4*���cS�P8��$3��x�o� �4�ro��B2�Kӟ����8�3ux{8M���߸v �/[�ֻOu�6����2����3O'���X)0�PM[�����3ȝ}k�%�i�$�+���X��zg�'���WTL&Iz�Κ�x��ڗZ���=U�!�%��ܽJ]��;KgW���v �!�؁���_�[��?�g�y��b�=B7�ҽ�N�C|���HY���=�c�奻����,4�Ȏ9!�;��%�0�Ѩ}��g�pU��:a�2�Z8�J^���ƃW��D�[|7�Wt��͵/Iٶ&�3��x��5-(�TJ{���k���*�콫�1:g�Ky'\�_<9�x
�h~���c�H�� �S����1����,":Xh�#�j@A_]�w�o�T��К��oP�>^���p_qx��'�c_7M*܃{��o�hjˮ�^��uB٥���T�Ӹ�PL�H�2�<�75!��i`�rn��[
)h[�<��&���~ߤ��_��=�pE� m�V��M�
(��@���:TPf�k�f�WwcrC�z���e_�3G{sѸ���H,ZO�fX�!M��J�+�3�ԃ(�F�ܢ��(�'K'΍�W�Le�c����u>!	��K6sZ��G�O�7��R�b6�1�wٳ��	X�6|dභ�6_��^h�-"+a�jt_g�����ՙJa�vL�N�>cE�J��3Ҕ䍝�,S��Ai=^���o��4g?ʣ����>F��J��3=��ĬxC��{�����(�k�ꠟ������`��ۿ�����J�ێ�w��%�%��L�U�S�7]��Z�E���zF뭺>�`�+Elھ�GH=�s���@]��t���<0�<5�#'5��;@�}S�!����7x�����')c� �x�t��g�?p	�J�wĆv.:a��#pp�W��5rN�������F��ģ�	i�ݧ,�����}�v��&��_�?���;�DƑ]��2��k3����]=$���G&�^S��p�鐌P�� ̂�[����`w92��U;?����6��(�ū�*c�j���s*��d"?)�wе���0a��#M�v��"A�Ѧ��:\�2;�Iɧ�e�dQA�(�(��\�חPP��c��ؕ����1\KۊwB���%4�׎�B�dW#��^Røf�o+C���ǋ�]��W��.G��� ��å��2����K[U�s�.�5���r���ѕ�~�����u�#�X��x�H_t=mώ��ۙ�߹�	�8<�]Iy,�ݺ*T ��<����F�ċ#.T�*S��oQ��U����/q9�lw�@=\�;àv�&�<�4�:�+��y�b]^]�V�(��m�zr�m�V��:J�s��e�j��s��ơ������v���
����%E^}8v�t��l� +P��F��->��L�����қ����/���=���*����z5�O.z�po|>�	�����Ƒ8�[Qww�]���A�	�{��	�w�m���V�N�3��&�O2�x�Ɏ;�c�7Ж}p&�4�՛i2 �rF���gͣ�y��Y��������oc/�+�``y�!n�8��Z��Z�T��A�w~c1d�*.+��,$�Q`�ZdL󂨢t�b�B�%��V3���{ϋ����dt�6��P��E�*�Sxb�\9@P8يv�`+�o���1��z���Jev�[���yDՒg��*<V�R|~9dr��=\",
�e51P�ިb�u��h~R����7	w�����>y�n�	��ޞ}a�^���)���𑺣�:�`�{���L2z_I�����R�`z5کЉ�C:������/��{��b؟�**�j��>D�=�����eԕ*lń�@�u�:���U��P-�Mc�!A�>?��7�
���:��o����Zbg()S)���{`�%��zR��Y�Fr?��c�~�̏y���K�ԟ�p?�sx�+����F|���X|s��x�dS���J|�`S���k���9�s\�`%E��~V��������<�K]��U�x�G�D�3�4Z�� �����,i�;������*��%¤�~�����K���T5@�ϛt��CRh����C���'��\��B/>�Q�)����3���ZKEA6-+�ϓ^���$�AK�r���R<b*��Ґ}+ �����{�`��MWM#]�6�֐���$����]�׈;)�ٛ�4���f���ƈ/��@�B��[4i������!S�C"@�a�:�IZ�����.������+�r�Q����i0���KN�S�T�I�xx�Z�� �b��af�D����X3��L~����D;
\V�J��X�~�`w��#+�7������.�X<��Hne�j�2��a���3^A>�s��ʥ�����c��;��y���q��ztxO�e/v�����Af�T׍�����J�.7�h�-<v`��=�O�R��EDA�w�IBt�g .\ϸ=Q�o�����8����x����K��eޥ|�a�i�s�HmC�v��3�n�ZZq�d0kx0�X�&��3��X���VΆ��3nX]6_�X ק/��'&eO�'�.N�)��6޾)�lT��3���Nq�[�Z�N���sH�ot�
�#���`'o��_;�Ҁ�漸�u4u�1��L��A��"Ȕ��;�t����|;=��"v���8"ɦ�7�Z#�����Pdhx�@�o��,�iC�S(g��چPc8�ظgr�Q������H�É};����
{�ii��hO5O����F���q1�e`�M��c|Z�J�m��~����p�n	���L8��� Qvݲ���$��3k*��|Ϥk#�7�̆d9V ��b��<&��l~�Īr� �I��d;U���#�.U}��a9*�`��K��b]��&�B���A6�)9��rI@F��a���] ��-�<sr����v�q��]���.V�<�ռ
�fN>��÷ԋnp���շ5�Ѭ�DF;DK��O��Q��S���2��+��D��F��N ��P%�����$9�K�KEC}��˦����A}�B��њ�1{A�f��݄m�J?pRd�
8P��B���υ���ta\��;A�y��ױ�{�h$��QQiA� m��#S�N)���D]
����1��c�F�r2=����_���$��;��X]Z�z�Ό!��=�ymt����v�V����~�(�:t*zp0	D;�}�J�A2�g�Q"\�+��*^�$�{XEh�*�����rYGԓ�
7�F�p�j����g�܎�:��������~P�Z�H}%9�c�?�f�gq�Gj�w:�Ȑ�_��A������Խ�u��n��``gr��9����Tٌ]]�f?#���h6L.$��'w�9�z0�o�HK�����bX6�,7(q�{����'nzS�=co� -���ԨN�Ϟ%�pC�e�f�Uegd�x[�Q�W
���@8?/�Z��h`��Az�~5���<	=��-�	|���Sl�4�K�v��im�>f<���;w����n�C{�)�*))���kh$1?�=�듓��c��� ִex:M�K�.u�b*�eV�T��	���¶D�l��=��%E`E��n�����{C�ed���5�6�%C�E"�i��Ӊk}��{+'V�_��g[sDV�����}
�ӱ�D�8	�4U
��FEsŁ�Šs��%���G�]�����G�l��c�z=�n�ş�l��yPQ&�D1軑��hI�Ht���U��@�K"�U%�x�ҕ]�.��B@��Ui��y�8C��!���JPf�y��	�2W@_y��W�!�I����I*�Q���c�]΅�e��n;i�2����2uj\g���7*d�	,S��쇱��UUxR� l*�A��(�Lsv�L����=3|xlexzK�Q�}!��_� �&vm]����AiVK��t�lQ2XF�Xk3Лt��P��<ﺗ�r����q�Q�������pP�)S,ГA ��!�[��^�iX3��`���A�"�R�6 ��q�P�}��a~t_-�_8h��_��
Z_ݴu�0�p�6��ҁ��՝�,{�puQ�ύܭ1�H���х�yD:��XvKH[���&<���(�1Z԰8̾�ـ�l.�v�ѭ�5cv�@��;�'K�q��u9^6��zu`��X f�_�����B���5f} Л&��O����J��]hKiPq��O,f��i]�C���t8%w�Vi�ƪĘ��{���=�3.P^S%�M ���#�P�����#G�F��� Þ;xa�l�=�؜�Y���;�/Y���+���GI���S�����7Ȇ�p
7�۰qw����o\A>)G�H���EP�<ʪi��.F� �9s5\.�*G����޺^uc��Okm�s��P� ��a�p�tV����ƙ3��!_�Fk��O��=��.����tθ�*�#GGT(�z|�.��#kR1�c��$�iw���G=R�*|s�4��bj<!/}L|ۼWa`#x4:VG���7��o�3�9����u�f��)��v
󳖗^k�w�|�O�8�V"Q z�l���Q�k���ߖ<[��N�o��A6�:ւy�#v�Ӥ���GQ$z�����a(T��`�̬�1�״�楝�7NI@%�8H�Q�-�0�k!.�GL���j켮��E���c9���
�f�?i\L���}�B�p`�c��a�R�F�{+���ݻ�<�n:$'�iP蕄
ϧQ?��uE��&o��h~O6}�a���'�"�8���ze�D��Z�k�����q��(�?����	ou`����O�q�ˑ��a���;���a�>Հ�P?��� ��ߍ� +�0�|�0
��v��RUğ�<�V���
2ɞjԸ��L*`�����2&��D)���m�=�?bn�ƺs�X�����FsH��~�����w����Y8$0;ð.jF�2�6�{-)�IM�������9ҁ�^��q��hu	�Yf��O�H�zCA�dteN��ty�&5�c�-.|T���}���E��z�ߜr�;dv�0)�6$�!@=�����l���)Nq�~vݠ���Ql#���p0ͼ);h�q��{S}7�l��6e����ၰm��L�1ܔyd���X��Ƣl�~D5z�<��M��|*�>�Y�0������`7�4�!E�}婱��8���/ݩ��ȉ�!�ӒH}=1��i��R��g��x�pI���/q���m����ߍa~"���`��|o�JxÖ茙W��L_%Jy����O� դ6��`�y\��˯�$���?��Et��ła�����ZZ�_������X^B�I������^�kw�@.��@��q�j�8;�r��#�Qg����̣#�ix���y���m���a��.���Z�I��3������P��7Wfb�2���7(��z��,��X@||�b��?���m0\1{1]C��'����k���n?,$6�*�w���q�ܳ�D~�p�/�6U���E��1��K΍
ix���O-hH%ݿܣ����D�S$��]����g�a������φ��墹�]Q��QR}�p���9�&z��nDy��+"U)#����l���ZMt�zY�>��~��McЁ
3S� �N쁰	��tr sX{�:��n8�J� �1D��1���ސk"�W۫?#&�$��eYq锌J��k7%��Fd2&h��AE��������=�>�|,��X���&x.��R'��Se�Xv��qf�J�:��.��k�$�B[
!����<��d�F�rZ�M�|��F��	��|�|�DZӦ�o�VA�~BV��J�p�A!���[�4���L�_����?<w�iň��9N��!o�&�Y�(�&fwUw�<#���Ȃ�C���vz`<~�}��d��U���_��1�ד$�t�@2�ZB������E$AR�ӷ�r۫���ebW�}u#��/�" y�D��&�df3C5)#������U�W$��
YV�E��֞��m�zhK�|;�Ѽ��z�!:%�.�IN��XN���
�`BEG�JHm�V[y_�5\���gn�����*�օ*�Ad�6����L���$�Ր���*�]����h)9��{�C3��?g��3bA�0���^+I�XG�!��B�tg|��`�8������]?M�2H�r����6?��T��߭/�$��&#9�l:�f�YI����PEU�&�Լ\N.%Ǌ��M��2(Q5UX_W��L��`�,�3EL3p[��E8a/l�i�W�;8C�C�P1{_.���m�c�^k�ԏ�z5�Ng"�6`��S�;�`�v�}0~�X򺶑�w�.c]=O@�t褼c��8"`-e�:�2z�}�!:3!��v�X��N��d��iw��j�Hp�{=�kG�4�Sk�?��B�_vW������C��]�C�	�7��%PCH�0wހ���|(� ���B!���a��7�(�.#3�DUZE��{�B���e��m�W5��CS�p���}�qZ�F\�)<�?_Z/O�P���iP�4�B�C7\���}�k�-�j�
W٢�<���;LD�j ��2��v#�p'�Yt�)����1M�]=����$�?���1j���:5|�/��J�J�7�߄-�^l+F}�ܭ��B�������Te�%T-KK޹�6v&Bch��G��ؿ��{���ˎ�	�\�dB7>�(O����I�dIx��x��� ����Z[&�6�n;���`1�����'��8S��N�DyM�Ȟ<y��e��%v�g��@�1�CY+7i$�ԭq����E�q�(����r�h���p�J��n=����3�sy�8,S�u|�栶AO>ws�V����Q��}9�a�f��L���AΠP��P�A�XaV��Dy������N��Ȝ9����z�%Y����#;c>7>��6@I��΍��I�:&lO#�V�\����ԴZ�熁�P��l�_�CB�i�з���xRU�]>��!=D��6R%樐�'�_S3!w�/Z�c�?��/T(���uf -�6�^����2�P��\�G7���|w�򷊅��:Ʈyo�O�]=�$K�f�JZ�:?>8[�\�py���n$�"L��\���hI�[i�\ 9#>�ϖT)Y��3ِ5 &��F^��@;uS�7�uX�->�.��}A�&�ݸJ[�҉�B�iұ��W�;;be��������[ȲY�?I�%��M��FZ����I�^�{K�#�k2��S�@y�nQzULxyc�ot�,Ȗ��}�mc���N�q��{jV|�J����q�w��J�3=�5�X�lMYw�zsbFeND4�la&�g�a�"AU�ؘr�B�_�݊���ŝ��#������=��ޝ��+/4�4�d�;��H� ӗ�D���)�JQ� ���[��ļ�j(W�Ѿ�E�4=D�ʑE9�F�!�d���c\�2���\Pz�_S�s��y��@�d� BT�'�,�)˱J��Bfn`���D1��Sf��?�|Z���/rJy@��2q8R�&��N�2�m��ScD�Z,��e�<(�#T��b>��cnY��G�yjJo�gjma�K���;�@
�`4���
b}
����J���Q����};��*�Id�"|L�`ad��5�Ke��ˀ�+�J��uI�w�Ei^��%�'?.��3de?l=0B?r���dp�|#�=�[$I0���?.\n���J*bO�G�ǻDcHൈ��_�H�Ly�4"�Z4�}�a�_`]a���#���s�A���|��v��Iqd=����`�lXE�B�cE+��ݚ����1����<��p���Y��\�s�-���OIBE�iRx��	@�w��-����X���#{���>(.媉�N��+C1��&0�y�0#�3�b����]f�m��!�Ƀ���$���y�������׮���"��w(y��|���ϣa���+x�۰"��5Mƥ���|�V*vL���t�]/�o{S��4�ĭ �=�}���=ѭq�.��%]o�����U���/nX�������Bu2N�Z�U}H���'k@g���m´����Q��I��E�]��O��76�sG��HEa�8~������6�({$��@<X�jr>_?ۆ@R"M�H�����N��dqs����\_��T����m@�����q�G�V̾�+�[n�����Yx
R2
��.Q���[�i�.U��2��]�Y�z�BV��Z�l�|T2�TL�eY3�`��ON�?�M�P|n�_�4�$��33�̑u�?[�����z!��ܮw]*}�%�x�P��ڴ	�J>��pY�������RA�BQ}Gk�b=����;�P�"��_�p�c�wm��k�&[�w�('Z��!���'�g_ 9�X�<=�W��ȃ��z?�F�Z����Y��<�P��)�>Y�cn/Ys�sX�C2N�B ��c��� �AT�9l�fT��z2O+�#�o�E^�Q�������}�xP��ԣ~K6�~�*�ԍO-=L����^s�DI�L�^Ȭ}��G:c�;�<]Q; z�������������TjZWҒ��7��H\2��H�o3�Dخ�7�("	�8�ע�]�2" oBʑ�kT=ռ� c�|�.�.̻�I�Xi�Έ\�&~{&�\��9n�D�x[��L��(�-hnڿ|O�5�ׄ|f�T1�~�6l�P��Bi�k�f��Q�.l����7��u!���jn$ӯ�X�z�ģG&��J�h{cTP����E�Et���SX���P���+ÀQ{��/�;��ra,�j|�vk�n}lz� �ZmA4𨨑i�Q1�:fY(`�G�j��2��^b��}��?�פ:�C�PC���
�~�L 4�F�2g1ʽ+V��'x���E*�PD`�t�3�;3����%%2�d��	Ø��Nr��|��jAw����3�?�\�˶?+����fTt
� �_�4�^W
��BD!H�Ճi�YTبJ���$�%����8��>�#~[Bc,�eҪe��
��Z�e1\^���z,1�:�b$"� I���|�1����>]��i������Y��2�6R��qV���.�`����u�_�W�_�r����U(G���i��LqmBXq�vI��٥ޫ�u����\����Ԉ��YAG�G�4P�(����8��ĆJԻ�"�#3�������W��Y-B�@�
-?�#�����I��"�t�pU)� U��#�e�Cag�6�'О߮(��PcM}��x���1�2L.��m2.1LK������섍P�
���,5��,��p��{\����O��}�|&=���B�%L�6�� f�t>�̧��64~����]ي$=��\��~{{R��$��vW����)1̦a �=Ì�@hڶz�L`٢4b���&�e��}����׺��e��8�1lű�
��٢e{�m�WA*7��Zq�Q�
b�@���V�M�H�ҎF�(-K�y��>���Sa���r�?�(:qh^��x �!+�N&<��ۃ���.��׽ Z3 >��4s�f6�׏\/��Z?����/��7�LZ���"2��K]-?A���Mh���Yz����OJ�����9m�s�sX���u���&����=�Xr��7Jsԡ���xmJ�s�rQe�K7 G=fPB:	�e��oi�dW&]����uD�^P#���#p����z���Q��X�Oǔ��i�g�+l�1�-��M"im��]1���	�I��<hH_�;k�����3��ܭm���4�l[�$"�[D΢�����imt��A�ugVV*ڝ�`[i&²��[Hg9�w�9o�ď���UY��
i}�tI���}���ww®�T��z������c��z��T��y��-h�w@Y�hn&(&ߖ��X��%� �`#��B�l�\�A-IB��%<���G!�v��cu��X�33��A���/��^$��X���v�(M�M��{7����I�u
���>)Y����.����e"�y�	>\�5���!H0+˿7k�elL��>�������e�z���c�7y����ql+��2�XHH���ؤ��;GH����Z�cgY�MI(�y��δ&����<8l�jZc���.�1���F���O�^�s.�:�N�gR��ۘ��"pC+�����W1!�W����.�Q����v�櫠8Κ��ڒ&\'�
C���H��G���&�	ؼ��F'Ow��,d�<����Ð��j�*ӭ*���ܹN<UA�T���Fk���Z9woH.�.ys(�g�]�I"�`�p�?3gbԠlհVhHr�)�q��6�w�A�B��n@O�s����֓J��/���آ!R�G��n�eF���=RE4�W�$�C�o�f��ua���s�N���1	g�� {�eW���ge2Z��t�hHoE<�9��H�J����z��1T�X��M\M������/[����0�6�E0Rp���*�lo�_5L�'D��s��Ac��~����~��$#K�7�1BXD??.vW�X�-�EKni-�Z*T7}�6v�wZ�������O��-4
@G�a�%�=���]xA���)0�f���^�7�rk��}����>��h�{ N_pu��'�:�^���G�d�]�sY�Yq�#q��V�����Ȋ�/����M��o�N�Z��ٲ��G�Oļ� | ]�6�V��V��Ӆ�.�sZ���V0�|��.7L5�K���a�W�G@�C��&��$pW���'��,���� U;�?½���γ�*����g0����������\��%�o��G8�/g��na�f��1YM��eRv�t�� �B���`r�X\�-��t0�җ�����i�K`�YoڕR
�]�8��ހS4aE#��Pi�ױ����l�Q���IS=��RC)_L�Z{����ncIᜥ�1u���Y�C���������F�J/%���T$���׿�2fY)�8�ֹxW�4k��nQ*�ܖ_�p��,Q4.e��Kq�����L�,3?�݅׫��BA��9j�0@���1�wm+�ù��^��1L�Lb���r�97�/�@m@�T��Q��-�g���_�ױ�������o�y� �pݫ]n)=��D�7~�O��I�y%�G��e��Q<i����<�a�-7��囥ߑ����N���#��V�6�1My(u��fC˸)��Y~p��V �9j�e� }
qh�b��[r�%(��,$��$�vi��ť���l��}���pZV<�ǒ+��-���NN�������J�;bjB�qP��q5��]�������'���-!�<]q4,���d�
�Q�HӔ��1�ֆ��E[c���S���.%=@JŭU�zO�6�����̊P�
Ҵܴnu�A����k���G��&��8Sh�k_r"�A��D�d���K�f�Fd��O.hG,��n�E��H)C􌀊~E%��Qxז��,�m�hH�T��x�����f�K������S��d�hm�\[�fQ�4���5��)
��?c�d�KȪm�f��Gt���e[��g\���s���{�xQ*]�MUJ}p�RҘ�Ʃ �~ i�kS�>�范�`�B,`�>���mG�}�A�U,�){Y����~m�_Fh���u=@Q~��&��u3ƒ@����!��6>�>���?���p����p�f}hY�d��릯���*;���+�%�E4Vl�׻}��i)YN��9M����x�芿�p��g�{d3b��,�m�Ǟ������q*��d�j+�ݾ΃4X���yI�_���E�hyA�B��0�Dg9�N������}�=�!,ؐXq,�7�T����㵥�mPN�
ό� s�PA�*�������(G1]!,�뻌���.@p�y��H��ƫA�����XL�4�>"����*�9�P酂��F�|6$k�L��o5��c��ҒVӄ6k^H��g$�	�8�z�"!=Bz�+�V!��I0�?��������C ��&�^� ����S�bc�uU2\{�V���gAe��.����&ŝ)��������ac6pp� �~w��Cߜ�9O���3��k�T*��|�W��"Q,:pTR=�P
4��#Ղx����ϕFi©����%8��9O���<9*�L�`6ZN%*��%=��F��-�}��Kp���R:x�g1�dS��rp� g;�"�؎񒎫�R�rUjp�oP�*�*��B�@�`��3Ą�а����!�������T��g]؅i�6w���V��ԃ0c/+\F��u��G"�1!��T��9�3��j�N|��{S����z�o:����أ6x�'�2��<0щ����R�-&@���F{{��*���{���;�P���������A䎭 I�{o��.w����M'_�	��g��:<�S�h��y� I&u��o=	�!կ�z���UQ��%=E�S5�d)�Eb~�����]�F��x0�@K/_���!3�g�`T7��XM��	[�Ӆ�y�b�cIF�qy 9���ɡ���{�?.���U9Vet�.���2AS�Y %é���{�Ĺ��A!%�^����R;B
�,8�,�,�N�)�?~��;F��(�\�A�C��z�V�z���zm܍��%I�.��U)nX���������]��!�X���z_�?oQ�%�����8P�G������w5?��V)�4�ۆA��7Y�s)f�ϑ.��3��������NF�e���|�J0��D�<y�c>n���٬��;�}o�N�[ly��L0�1�g2ɦUp����x���n���	&mEP��IS�ځ���%��O�H��X�T��3�_������� �e������-LJ
��.���l���g:�ې^j�p���A�?�,n��&#�`�|�w_�v�;{2������Z',���Ό$q��`��n'���CFj��(��8�:����Wwv�3g��ڀ
�����56�7�K6Q�~5h�}�{����Y��!o��MTx]f��	?���ͅ�\T1�<5Hr�%��}٪ό�d�"�\-ʩ��r�1���n���/�5i���$�^Z�U$o�Ӥc�P�Q����{�dď���ā^q^1��"��WCW��2B��1�xM��5���eJ��/�O���D{Jׯ9�X�Z���WK!?�����^EH��\'��/�۵r��Tu��Cē�͞��X��C4�0Ku��!g^&2��|8!J�ϔ�E��-wo���!*�%��3; �&�F��M<���m\��U�H��jŲ:>C��I@"O䍗=�쥒�mU-̗�T�����d�y���@�VX�P�:�@��YfêM��1� a�n�L�?�Ͳ��	�'��v��c��zGr���ۦ��HBe� �Ť~��H�e!.�\�b�s�1�~^��0��c����C��H~^�
���g�swm�������ޠY�=M�g@�n�M�6��	�� ������h�|���_�l}0�G����'�C���K�5���Td�>��'��{�
}��@���ljA�R��PAeX�4®l�9����F�݌0�\�M!��#0M�,���Wg$]��ǆ�~S��=�@i6��o%!ۀ�P��_S���Ì�pf�b�&��� ��=�x̅)0wlo�=0��~��v1x��5��0��#��X��� Щ8�sB|O�gpf�#��ؽ�(����~yT���f�=oCΕQ!]�f�<��U�ae4Z�f�Z���n���U�.hKC����H8�H���Z�������vjv�-�U��@���.�{�,mw��DԹ$|�󡈹ֽ �4aR�����j�#a��@�b���H��PB��K%E9;���k���|�u&����wM�R`�Y��\��KK�L��V��KYw�s�s�n��&�/H�m���c�R��B�.�1���>�6�+E^��IBY/n�˘�M�4O;J��m���! YݱdlS��L�킟�V���%��픐a�9�)x�؏L��(�n�	���)U=p��@ӹ:��c~���Xb����jN�������m��H�-*��n͡r! ,͈r ��?҈`Ůz�_b���;��k��Z菅[�Y�acTVj����M�I��+�D4	����L�NȢ��3�º�6o?�z2��Z��	�^in�]�D��z�l�� �P 1{�4�Y1�<�(ur���b?��G���V9i�_��ي�F�7jQ�'T6��'������%�Rz�ȃ�w�ˊN�����+[P^S%�Kء�Gj`(�m'%E-��$�M�p��2n}!J�`�7�ǖc�%J�=5g~e/���/(]ְ%�FEyޝ_�zg������cv𢹋Ɏ��}F������2�GEz+d�:{~�q~�[X�}��V�9+�ܯ"��8:��-�s���3���"��aop�yˁ�V�� � �tIX��1h\7�a������C!�Ŀ�/H������z`�?�Y�L1���\P1G�p� 	�_jJG��<P1.��u�{b���Z�V�C_�w������zZ"�)?���q�x@l��8$Bz�^�5���l����1���W�\q������(���-(X|t�e_c|\$�8f�ov]G�f6�FpI���I0�I�/8�b	^I�U�*����W9@I�#ZD��8�E���&I�,�
Y�	��~�`,�H̀_��ً",�e��|���P�gW�2�/�ީ��H0��|�,�q*��z�t��Un/* G�:�v�u���s����)��,!v�Pm�FzB:r��X��aFW�e�S|Ħ.�Y�{��ͮo�t��<_A���� �Xց�{��O�%l t?�E�yb�%nGV}�d�_9Xg�v#�Le񦩸ޖM�-"�M���wĪA@c/K��C������+��v���@�.������̈i�9��
iFË1���E��/ߢZR�?��� 2<9�lM'�,��6��-[�0�d�&"5�����E*U��S�Wo�V��x�e^!�<l�/��{>:�c����c=�
B-j��m�n8u��sE�J�]���mBي�y74U��+˿H�N.��S=����c���/��u��L���XYl�q���.�	!��(C���[>ƚ��j�H�ř��,�Y����h��:��IO���L�#�а{��g�ɵ��S�/(���gd��g`��f�qçayx�vj;��>�7�d,ɱ����H�Цj�GJ����x&��~[��p���I�h�#9�SxB����5Ҿ�b���7$-�CE_������CD����i+fX�W���g��E����Ini��}FӾ���}��Vo>�8$�����!�ͫ����A�C�mk�9ҏ��.'aq��X2�};}�ԫ$�TΦ߂�dCnO�{��*��`�z]��	o=��9��ͧOЂ/a<�DS�L��^"İ�y��q��7�S~������^=�
��V�eƪ�y�5���i+��i�X����Ԟ��@����Ⱦ����n�s�|J��K�����G���ژ��	��0���'���<L�C�m�5=��K���i!����)������	2d���uL�ο浿I��B� �(#��^w�b�:+����&W�U�+��#*�U�DD���+������h)�W�΃2��y�1�	�z�}�����6�Ҿ!Yr;Q�����\q�����^�]y3�ڐ���&��3�xk�6a�,)j)�y�.&���Ux�#��O���g��V��"6��`��������#G�����q��m��r.�@�X��f ��:���P>��V��^d;�z%�ۘ�J���@$%�9g��@|��J�M�xGL^��>�N�ԍ�m`�`D�cd~�J(�.xr�k�{!�܉�$�'�៉L��ҐN��	B�x[��O��/����Ʊ[;�EK�ٻ��LU�D.ߔ�R�js���[���9L�x�~��7�N�7`8����I��i�P�YSg񨲤ڄ��Na��t��;��'%)>k�!�	W]Z78�)
R�y�,��y����\{�䚮��u�
<��ŲW���
R\�8��U&�
�,��X&���W�_0�su߫eO��+hfl%[I�����(�<Y:=	��D���������^���.G����w�o��R�%��?�Dd�Z�Dz��w����-���[gBe��+�IG��-�<�f�S�s)�뮞2�7�q)+k�eX�O	�haRZvR��A�s�J�i֯e,�z�WФ��~Fr��@ k��pYzĚ�ߞ顆X��
R'�F����oG1�/t�B�b��v�ކ��ё�Z�~����BO��𢀼|�Jl̑�{�E�%�H��驫T h6��D!l��XqUoКhi��
���dqz���m��:��*��'_��C0��a�H5�MwPL����"S�p�dX�x����L[O��Y*�>��DI���_�{?�X'�N�K^K}_�����} ���eETw
Ij�j[R�Gr�dS���)�Y�y����O�w�/��=�M�
�/�Es`�pH��{CF�a3ї�O�ƻzҁg���a3�$FZ�b
fǍG����.�u73���Yj⯢�g�48U�g��ťX��!�hݛ�p#'��vWзu���o��;�J�s���L@3i�{��}�N�xw8�M����b:��9v��o7��2�V��h�$%VD��`k�1���A�O􊾯S���`��iW��� B1�������D�fۋm���{��x�l��DK��H�*B���ǩ�� �+e�e6����{�&��!�	i5f�{�@{�!"*j��� Sb#1�S�rP���ua���?Eڕ
�.���q ЯШXG"U��|~*��x5qP~p�U�v�V�z�?�������=�󽜬UY��A�k��wҍe�$�Yo��PXn��w���6J �`U��A�E�����p���f�7hy�����E�|�	��3=E�.�,B�����x
�F�*		B\�$���7�	p� ���Ǯ in���E�u��p]����
Z�G|�?�b�XT��'��:7=�'[{>�*u��*Ahʤ�&�ε��	�W.������� ��2�f�0�&����Afh�1H���D�b��#(����=F�<� (�i���Ռ��,�<�pj���#����"h�lp�]��4,9;C�@<1��`.����	�������{Ȁ�����5��s��H"$+G�'�D�ʜ�h�Y
𠞱�N
�z�B��>wUX��N��ϮлL6�����ƻke�t=>�O�:����P'���~b�C�4t�� u�����\$���Na�Ҕ���{D���
~n��ԉMj�0&�!cOWAo�B��KBl#�a�ʠ�����{A[�!��p5I���;I�7bY�=&�M��D��ǭ��'a��2����	@�t��ѓZ1�#�~�L�����	@��0I�������]�����R "3�'��ǿțf���n��B bdDb1U[������eR'��dhf��k%�z7�g�;��D�Yg�E̬j҈�MxB�qE#�$'��Q����b�L]MW��v�=��zN�q[Ӑ���K��f�ro���r�ڙ�L|~7�
���_x��_�C6����'���U/�y���쳎M�/랕��! m�b=�6��~��ٻֱBə��KN�[��2�+J2z��8��������&Q�}�(A��8ve��:6M�6%`
��<2&x��%��[V@��M����,�I D~��&�Yh� Q�ԙ�5dglߴ��E�O1�����=��M�];���0�j1��3�z��sM�sm�^� �j�#&�+�W4a��������ox��۬o�~�#]�hE���#ր���LPUIz#����.�����o�4�O�n����{<���K���3��ެ�3G�2�߳rI׹[�s�ލǋ=r�9&#�~�;�����Yiǆ��ݩd'��r����_f�O�m
�Q��7��KU�����A$���\&8��.�&:��T��v��@Ka�H�Ib&#��)$�v�"��	+>I���ɚ�Yш�MI/Y�!l�̪V�g*m�[d~� ��
lp>�7$Mn]|�$x�����'���J0-7�FK������5#�#��ňc�p/'���R�Yi]`|ǒH˔;D�-@����&�) ��s���8앎,(EV�� '���̤��o�4h�.�8r^�����	�D�B�l*zd���b㾤��s�������@Ч?�P���AMd��o>��`	�K�H���S�&w9|��︕�J����;����a
]3��SQi�G2���+�=��v�����Q�����L�,���kUp�e�+���U
���!A�/�	�qG��Q�B�������F�q�iĉ��N���S�<Pt��8M�^0SJKe�'�8��%
�5�tL����W�r�p޺>d��c�<¥fK�\Z��R78������/e����3�K�<�����f��ߡъ��Y.�RA��&ȭ๮U[)X]�ZO,�gU���V� �۫= �9��9FGZSG�`<Of�;��Z�{EP���8@�Oi����o�'�K����l+�E�E�?`� �R�oJ>��Yۉ0��:i� �l�ُ����-w�*-�`E��0�/}&��n�B���	�(�K�u/���ˑ���ڽ���q����/~R�g���Ĩ������n��=6�f.���ma��QV�Ɠ�q��U/Y�+k�X�%���aK��r�4{��ּ�9x�#x���|��)�tOF,�hF�Zm&�ۓP)a��e"�4|I/�W��e�)u��@f��.�P�AILr��`	ap��H�]G<���6V+-�V�푠����y��m*�]�_�;I�7b��W�¼+�=?1hE5[�u��ܑ~	P�P�43�+�˧wd~����Y;z`o#��8X؄`���|,�G�V�KX�?~3*m�(����\8P�a�l�U��R=C
���
�v�3m����gM���۝�Һ~��بW�W'q�svW4��1��Sʗ{5S+;F4�K��������!?�(,� �s���-ch�'vC�Sj��oJM�ĎƟ[]�S�2;�R�6�������-څr7�A����v����DX?��b��B��ck��zK� ��G��� ��ݲq�G�뀾��3E������oQ)`��|wLN#���V�d�I������וּ��5�Gn�S���z�&�)>?�po���H�7'�"g���y*���V���?��y�w�%2$�z=؛O��u�9uR�xV�%l��ƅBD�6^Y�Gw��W�V)v����ZA�Nچ{���	 ����h�� Vfv���݀�^��^ףH�&*� <��9�M��t�x��2ů'"2��w>P+�h/��v۩!�-�ǭA{�qg�<i�� 
٩�u�HW�%ԩ~,	�O�8�9a�ZC�� ������-���p�-b�3Geyz��𿟖��ָ��tZ��z�:2f��e2#�1}/�%�S� ��qI.}��?�E��b��}��3	�1ך���Kw��?�C�p�z9����ʟ�1�w�|�*)�bGBU��]u~���)J8�>)��)��n+���+ ���.Kk�N��
���kH�М��������<�W����0$����� UH'����0�R{��S��6��Ž����[r�;�ck�&�ʲ��Ql�~����ճ��$!�ew���$�r��>�#tz S�*N2s�Z���+�?! 2��:�,a[&�K��3׹��f'��g~M�W|��u c�4�?�n:���f���fԙ�/�� x�Ѵ/���uI�=��k�X�;/�]��;g���\��)�o���Z��>߶���;G�0�V�ԓE]	&�Ǒ�%��Uc�~q�P�=.N������ƵF��\ݣe\�_s49�r�I�]�h�A�~�R�yX�;�&ԡk_u
3�=$\�x ��ÀFq<t(�'UK!�z��q.?Q��oO�q5їd�I�rV/�c��ĕ���5);��@�ms9>L����S*L~)�M$fÍ/ZM�v�d)=O_�h?eߡy�dmE VZ�ˁzG�3�@�W_�!&���Uղc���[E7��j�$rA�8Gޞ����R�3�*��1��s�ި
BuEO��o�ω���<�2!�T��ذS}�� �f�YB�%{����g������|�(�?��`OR�Pk �>F�F͂���0�[���T�w�Ѝ)g�qY\��@.���@c���*(TLۖ���n�	yI�-^��d>��P��|T*lu餹���1��"��դ����#M�^),�QG ��d5�0Ov���L0��w�a��	�b�D�
�qc�6�~0��3tf����ǟF�I�ؘLi�1Ť"�2��5��k�<y��5��ƫ��^���8�#{4$��S�bLh����>l��{���4i��^��RM�����Ϳv�*����4H�dDT��Wm�R��^����c�"�$�:�.�pM�k-�[��v�pS^���6��
������o����/��(�U�m����m�U��� ��aũT�ӋA�J#>��*��剈���j�P�-��/�]N��x��p!Z��U=�[:������(�O��9Ƣe�>�s��O˗|�=�3�"����X�^�@J�_�P%L*�4c ����&��t���
M��}@���ʹ��Z���`�X�\����;,7�H�	�Y�|�d-��H��t�u���Qp���)�7$D~B��V�m�{�ʖ��Z��=*�M�Ƴ1:���6��0*�B,gl2���%A۽�r>��kt����n#�`�}�U]�q���\��>�ɱ0�J�Gy^S���*�-&ɨ�db�����p�JJ�?���K8�7^�F	^�!�?8��Hcc@w�j��2�nlJ6=|p����(è1��F!	�P�3�t(��ێC~�I&� rJ��H�/�0�}�0y^���9�(z�}���sY/�"j̰	#'�52�6>ՎZ�:U�>��3[S�.�9�u��A��yy�`;V��Δ��g��v{+h��;	�H�}H��:��:׋�[k��>"ֳ�:�e��<^6%�z���FL�Q��:,�>ߨ��&�!X�� J��dJ��U'�:��ɚI�����|���EN��}A�z�C�\K~����������<Ns�R�I�oj�;�D���n/p��z�\�Z�:����>}˃L���}�x��=1��S9�m��j	�=^��Xz�ߕ�p�J�x��\�])��c8L��#N-�����8��雭i�cGvIq��#Rp��m������)F/�V�L�y��<y,i��Bh��a��qwBӝ	��x���6�E��t$�I��ݑK�����	�m
qaB�f��|���}�ˡ@��Go��,�Ɔ����9��xnC���&���:	59H�A��Q㵙(y;���`%��Z�Y�p�a#R����:�o���4���y��Z�K�������3�S�����ų"1a�"�������}���Ͳ����C1�ٲH�/{�1���"4��00Q��n���J��З�K����`�[Vi�*��t�l�$t�i���(V?�����Ŭ�f3�I���+1�%5t�׃���zHĬ���Bj�Nbߴ���������r�XU�'G��qI���ʳ��=B"h&��������ʲ��⧵�����Y����L0�2A��xN��)�(w)\�gW�ta��7 3l��"D���H�:dɳ��T��H����!M�����qdb���J�=qar�����F&TP�<����49D�L*8������M�pa�;�p���q �B���}T�o?nA�Ϧʚ}�����������m|A	��&�;����kN�6&-�ltԞ�M�ͽf�6�MP�:_64�5�a�B⦚1� �jڠ�K�^a�,6���19��)7o����)	�:O�6Cf���#�ya�3���fAp���

'�!����\|�e�_�������CMe'��Cw���x��!�5[A��v�������FN����Hy�j�v:hu�B8�i�e�����EOk٧&�㾰�S� ���9�f|�f�N�����*jBM���/rN���[�?I�5�����<�M.[�WV�%k���Ųa0������H��ژ��H��m,�Ut��d}6�2)}�/�p#ez;�����R��>:���`���'��m	8�|��#H[�K��Ἑ�Dӹ�i��#�ЃC���8O�\s�֟�/CӴ�ƞl:���}y�La��s��?��g��%JQ�f�QA�ޫ@���ިjF5�A��j���=Jl���N�;;�0T�˦�.Q0ݬis4�X�^c��` ��U������i�b	�I>�{V�,�!lQ.����<����Vp��mhsʮ���b��w= ���;z���0��z�@���'�DԻ�<��)o�[H*܈�G���>>�[�X+���JC4����@���E'����qe��q���wt��M���ʉ�V���]�J� �J(�Qn���WU�e�K�/�*�w�����2�7(8�i�
CA�SU%m&���4�|�G��l+=��;q�)�D�F���H�J<%ٴ������~'!�QU�!1�3�X�O��'�w�7i�/l!���l��͉u�2��&J�J1,m��@�#������������]p����}����|��¸t��]6��Mh�-�y(�}`�ȅ���n|�3eYK��q�ﺦ,�Qs�ki��.�4�!o��Z���{��B�@���q�������-! �çtA;Z���H�+/��3���][���Y���)Y��^#c2[z��eH�ٯH ����FP�#��ϸ��_��?��dS����kD�y�I�\�t��3�jY��}k$_�Iσ���? s[�Mc�/�ؚ���L����T�𮏢u�8����t���a��숎?��� ����/4t0��8�c���Z�
��x`��|��g2���"�Da��I�C&K��LY�������T���4���l2����qA�DFE�!�$��:Y��$�C˵�'��_���rTk��{��ůJ?�t�ÛfI@L[�Mv��}:��/!��*�B}�M$~U��گrNY��M��|�Y�.dA������>hFF��E�+ k4&}eEs9y=RCI J2��([\��	�?$��x�t�_ț��i���j�O6�^5��ʏ�P;]`"o
�RDx��'s��dc3�]d�M�Y��@��,W�:S�/�__���1 }��{��oG��?0n��6/K�2��q2l#-�������_&�V/s�q��Wu��p��b�K�mBQsj ����#�~ػw�~mT̷��>�K���C�9�V�%����D*S�� )A�+	��	���L���S�BŁ�t�	�
���Æ]�~:�I�I�a+��;�ɱF ��~0���[o{GO�9���GZ�;�/-����	�eX�<��?�|&fv�S�A+%�S<�?�9������X�j!�v�/�$P�2#��dRwV���e���@���)U�ƬhS/�U ��ߞ$���ȱb�S��{$
�k�]Swm�gt쿓�e�_��ϩ����Mz��f (n���i�m��ڂJx��.7�f�� v��TEO��AbR���Q Y�J�N#�'�c��"��D`yWކ���	7��Wd��TFU�w��r_�`Q.�ʎ]7hk<�j�|0O�jED�Cm��h!��d�I�G���dG��Ѭ��=B����x[Ъ&�s�w��KR/�8��BV�vɚd����$�U�~�Ԙ�Ŝ(�����)0+��n�[�r޴�2:����Y�����VU,a�.Ą@k}w��(��
:�Zf�\w�� � �����P :G�ЫBOB�����bd��WV�]�D�雅tn~�}�[�ۛ�+-�"�1M��W\��&xG���D�T�4Vv4���2I���[3;�-�m�� WY���36-jq
���G!�x�:�����A���e�E�\��A�طp���9!���Ӏ�@1�x�Hlz��Uy-�F�O�����(�߄�	���4i%k ���;S&�}>L��K��G���M�H}�rL�.q��T�-��id靡��-�	�j����X����#o�GZ��S:�R��`��~����Z�+�>j��?�;8�Mn�n�5?н,���EͿe>+��jV)�Q� 9+l�.tr ��`���4���P^V�TB���`�o����t������p,��4�����o5�/�7���t�Q�3��x����V<xR1%@��l��1P��4�H��xZ������q`#�Di�l�,@�g�#��F��i�II�G�b�Yd����591�̱2��� �$B,MHM����0U�Sm���j9�ց4�}z�Q��������������sC�D��&TjE�^�i!�I�Jl :
U���T�#�F�Krr3!�sN3��{.K$��LNMa�"=�u�C���p ����O�י7� �\�F�! d�;��])��/�����=#�1�u��|�0�mY�[�#^�gw�翸�&x���	J�����|Oq	�m��{���e�;Wd�c񣾠�;D;`8��lVa%D�n+몂��//>i�@w����DY��&a�9C�0?�.��g�[�P7�iZ��]��j��=m��i�����*�~�`,~��g6�˨yFI+O��3a˨�m�@Dɸc�^�'�^4�Y�;z���Y57Hm� ���x����pC0�c��Q�ǐtǮw��>�pR ��Y��5��1*U[ow��xέ��"0��nHb�����]Mr#E��载��ؔ�ǐg�V��6Gg+2�bW3t�S�KD��_�Eu+/�T�Fj lf-����	BBÃ���b�v{+�����<j����ؘ�xT���h�N��5�G����v�\���b�8Xd��1��(��V��x^��6���߁�탷�:-F'��G��KT�����P�PF�y�d`^���	�C�Y�{���׹"�*DԦ��ٰ��"@>��.I�>�M��[�-�|� !#�`�5P$�ޛ{�'+�V�[��V�����b�ϖڢܥ�{��<�D��B1{"+&����Jnȸ.�G����H<��βn���\�F6)n*R��9��Y2'����iÔ[8BM�Yg�e~�ѭm�����{(!1}j�8s�r�2�Áy�l]a�6W�~�5�D��:9?��XE��X�HDATj"}�+x0�����>�V�N�t������H�Y;f�V����H\�2�utc����&bN��"4"kF�\T��������n>MhZ��3��\l,����~`B��z-h�{3����r�C��צ62"��j�\��ų+�o',�/tm���V��D`�����kpm�۵�䴷����r��2M�������VQ`\$�m�<�:B�D�
�⽄���32#H �_h޾��|���SM��4�H����@;=�\~��Ø`HK|����͆����sP~��,�Gw����'��t�I�A�4Y^;�̀kBb_q�V�a>̳͊+~���>�HM1��_gw�& ��-��N� ;'�Ur��ST�|��+2����}�B���H� s70$��`,�+�.�
����j�6��=޲����=��:S�s��Be�N�.-Bu�����2��������T>��/e�-��w�(���Wo�p	1Cw���p�H��X��-��rN���&_���*�7��}Ց��[�+@�al�/
��������ʘ;��̕�aql{s�p��+��5�_J��$�T�R��ߑdg곟H��dhC�����k�
�e�2O8s8�AB�3�M�o���+�SU6�fk�[5��]}>ai�܉����i���ʘ���g�U�X6�k�~�ݨ��T2ʏ��k�
iy ��J;�+�_2Z��n� ��I�4P�dHd�~A�sJ�*Y j�O):�OwԠ���щt�Q,F]��y��|���d��b@���s[OK7E˜4���^��p���,���+k
+�ݶ�4�^�h�O^׎,�h��˩�&�����u�z��K]����^�;��˝�uR<$f�5hȤ�_�����f�4hKADF��$�J���$�/�4�Ϫ�2tгmH-;��i1o_OC���@ʹ*���釚��i�D�Q	��]f�M�pk�7�	w�d���M��Ğ$a�����b��+'����٪�Ē�;��>d��š־���N�;`�֬�M�D�	yۊo�i�����2�('d��K����9z���7�|���D*0&W{������.�$�S��C]=�$��ņ�O2��L�3P9��׌��q�v[�'[�4Υ:�ݐ��S\P�ϯ)}�) �}�ڒ��L9�������>�J�r�T�~��cqat���Ԑ�`�ͦ�ӎ��>����������Yo͸1s4��7��^(� �F�^��=m2�z��_O�=!C@�1K��9znĎ�{$%&�[��%Y볽�[ka,�6p�=*T���FR��kQ��}�a�CHF�+"$����K �аs����v�эC���4M�C1����zfW.��NUވ}t-G։f+�q!89��VUs��5K�++
ȫ����S�'�N���}{8�ԟV����R7�K��5�]��WB�w�k���:�]%n�Ԅa��L���M(4ei�U�d�I�� +�ܟ�Q ���=���\�7���Η��W�d�P�n�O�(CTw��-��U��� P�}W��V��.���4b���ұ<s�����V_"�qUL��ZI��#�P-I���:��C�h��!�*~�̛��=Ư�dﹽ��1�	q	�?�P�p��-�b��]G�V �T�pp|��3@�^��Ɲ;�b�J��,��L� �Au���v�� ���X_D+�*r93+����`5'�_�d/��{(2��=g��W�7Mc��1J6ZOɕ�f���:)���6G�kTr�p&+�`4j��Gw�J��2�NR���4�u�����\�����Fް�&������g��>�D�}9��a��Ƈ>NY�$�2GA�+u���f��\��ؾ�.�-�G3_���J
����iIӘ�n�O�d�R�I?Z�ak����^���<@.�J'���:.�Hc��x��!زܓ�.b�����!7���9�)q�O-9.c�q6���@o/$}�&l���1Θz��B��'����`%}��gS����ăx����^��:�:pHq{�'�|q�b���n��"����K��ȼ)���9�x�<P��v��\Si���O?mҰp0�?t����ح~���_[g>�\[0�-�U���$�7�ؤ�F��Ta`nm�L��F���N�ݎm��.P�����:�z{�2�R}��|�용�qR��,�;)z�e5��|)v�#��
0�i)_N 8��	�XMa*���ڜ���a�N�������\����:�4?�`,��C���s�l���Sָ?�L��<)�&|:G�)�pl�g3�;Jy���)����t���{wX#V�" 
�d�R�	G���b���#�i;w�7�U �& wp���Z�{X�T��|"�9�Hra�x��'��U�_�ы���YP׵H�K{-�\8��䤨��ߣ����I�-0�&�֙b�5q
���gF��� H��
��]c'�c���ƺ XE�����L�~�������=�f���I*sM��/�I�����*�.�3wj̄1�Ț�['�Z�[�@N��N�?�89�G{E�(� 	^��{tw���
�k��q��̾ʛ�}��6 ��lF��g��($~�E���TJ"<327�?��� ��E��`��a��3�~��*"Ci郘�z[$nܑL=Ej���]�N$�k��,�pQ�!GF����&�&�#��Ե.0�	2x�ɡ/(D��%vP�f�ʯ��# <[޾�yU�8 ����A)���cF��V�gU�Q�(����0�  
��-�ς�B�}��!����*��)[ޗ����_���~X=��V6��,��U��m�G}`�/�m�BS�r�17J%
ϳ����vq3!+PV�w̟��_p�ǲ�� �RH=C�_����=P����j;Xw�Aj��rU(��}��'�4_1��̳H4�'RM�_2���-<���8�}}�	/S������H���>�
�3:�)+}�T�Kyƴ��ҩ*~��OM7���OC�`W�����t�Ԩ��.S�$�e�N�WK��8!�R>q~�f%`K�V�"/I��,k_�oT�*�95;ܘ��W���vv`���x�y�E�=��ԓS��Jc���5L����$�=�4\���uo�����J/�h��5����!A��:�o��J+&�&y<�P�	hI	6v�Q¬��(J�Q�wI�l���Qk0o?�:�r�2z��֢�^>/��.���0�ӥ7��i=�j��6�t���'�K�9��N��9�񛩿a��YmS�[�W�.�@�R����)K���9�G[E����&��2�#)���"hu�-c�~��t�hP�|�C�{�@]��W�GwT��2�����ٲ�m~$�����w@;&�ON�i<#,��+�ec���ֺǆ�R���?E&���z6�6�6��z*��l_�m��qQv2�a���aq�^���b��'�A�N���D���I�����J�>��]��?�v�����bK�
�'44G�OzR���U=ǯ2I�?����R�B��+�Q��E�m=��{���/����{��9���Ύ ��*0}h�`���lo~�V�y�t����#q]mH�0=���HF~p�N�COA����:b �9J�1v�ǁ�L��" ������1_��Ī�0b,�f^��8xf�$qh���υY�Ej�l:�)`P�E_v��
��-�G���9�a׋�༥p���}Hg�F���1Is�DL��`6�_����VG���Q�X�^l���J��ŝ!�EU�t���!����s�B1���I�&3?;�9���2B����`�w|p�-�%³�3F���!�}���ʠ�;�ѹr@'.���W
(���<�e'D�̉�p|> �M0��q���� }�,]�$��EJ��!I8d#D�G��J�n��mI�5-3������[�)����4�k���fM���-�c/�ޯ6�1ӿ�EЖ�FwAj� ]^ˉ*-�d#��j�8��Ħ�+�y�t��dj6|��>� �v2<tb���u&�60�Ga��e�U�2ܙ��[�������Z��zM�MQ��S�:��#S0tc@"Q���1�*z��Wѥ��Ƿ_�q�x4+�.�Mp�s%�󊧛���.e���Tw��iP�IM��E��D���q:��!���$"�������)���\/�N^�j��!: L��8����H3"��u՛����b�~��uzoCU�u��C
�;�-�#l�����m�ؔD/��4�_>6��̄5ǿ�?J17���{�܏�
2���\�q}V߉:�9�D���Pq�>T�h+�I�`D�F#� �hw�~{����N¤�������3۝`�?�zvt�T��]/̭ 3������ö�V�ID����ι�3u�2��W\�-�7��2���q/ u���3%����ՙŶ��FPR�Z>��*��SC�c����
�����Vc���\�R�{��I	�#>L����\��m{�;�:�|�h�Y�x>)*���m#��[o�� ��e�T��p�!��M��8�ls��������C0-Dn�8�@/:�@#αÝD���/�ߩ-�\>Uv]����<C�u���X.'.���$�JK�9���#����ƛ�������q4�n�9��"�MI��r�t~(J
�+U,eKџ=F�ސ����a�߹e.�p�>S7��Y�冖�H�z,T*�0k?恢ߺB�w�i޼���`�Q�E�#ow��]�ec�%Y�W`;$(�jd�Bhb�GJ�rP�K�y^��~k��c�ƥ�Z��B���;rpB�?�|��;w���V�I%�LIC����^n݉y�>(�9� x�6���a����5�k�T�/l�_�tvZ\r�PPO
THB�w���c��y>2$/BnOX�zj;�O�K����zR#�����;�&�4:���`
_)(�j7��HLI���1deP�ӐUw�s��.�P��U
���4aS��ra��N#99��@�6J%ׇ�WM����w�c���,�ᓛ� `KR��w��}�͔���F��I�k�|��2;���A��]�pPn���tCy\v��\������ֽ"�9S���!�U�Bl�fqѺ-\�s)e�:߅{��5�m»�!w�t�N�Ԋ��3�?�p�F#�R���+�5E�W�+�7��x	�A�X�����=��dB��1B�TlX>����q�.�O���z�BߋO��Sq�}�`v~�u��.�{4�d*&�'˫��Sm��8�� *�~��W�e��F�@���zo��օQS���i=�6��K�v�����qRO��7�q-�v6Ȱ|���|�/�>���%.���ɧ
���c����4��ԗ-`��9���Q��X���A����:D����1�ZX�(����`1V�k�GE����0{��Db�ľ�1����P:��ӏ����f֮�����3ȿ6>#�ʖ!�\C��+�������z"L=�E��季�]SVd�4��Ei�V�:�۫��R�?����"����\�?	�l�� <����L�'N���Nd],Ԅ��>1k�Ә-��e�9��|�k��>S��^�p���Vl�n�79{r`�?R%*x!\j�m�,6vV��˶+��U���vشY���Y�w$}S�LXN)�����p��|�7���v���|`�i�V��9�X�if�d`����܊��&�ᾮ�V�z��J~P�/��
y܋Xz�N�I`ͫ%���|�_�� �y+��Q)�;�阸g6Kb��2�mX�o�+����$��VSwR�����+�������^����x�iUH]ώ�{m�6��!��͆��B��ngY�k|���9&-$�&�Wl!�e\qjC�a��:rTD�������ɐ�ˇ8Էu|�R��[���j]�N���Mbg�`�f@��GF|7����q�T*b4�Y�Ԁa}��p��=��}1�QU�"ӯ���M���C��=����I����26�b�
�����ivt5J��uX�g��ց�|:l퐃O�,�Q�2e����}q%���4� ��������v�o��lt�!����a�6��x@6"���+P��aW?�0Q�l�JM2�%�J@Ŗ��m��(cP���9��2�s����wcs�B�7�Ѥ�'��e�7Ɵ�I����:�޼�Mr�_���|��"���c�W8�fFz\5�b�>c^�/��9Z��<��<^�]|=gH�3޺��<�)n�^ڽ%�A�P
!`�\Ng*�N��R2�� �y���aTuHҧ��j����f	E}Uҷ�Եr�E���\��N�ŮH�M�B0�ȃG��YԽP�A�����9�)�@�>��-�,�~�~��!s�a�޽��\��B��׳��f%=-��k��	��x����eO��WV��i���^��������b�u,6a%u���hHVm���49'Uޕ�nWL*�j�Z��՜�/
*��C�Иpa�e}���m=h�y�)�ڊM�%v<��g(���ت> Ν�%����uS�|O�\�� �~lm^Z9�VU .q�)�r">��+B[�����YS�!��/��q���-����oU�^��v���s�{�P��8��������3�9��y�sn�[��ӗ�,�#v�����).���E���&R��0m<��W����r"�sƀ1mEs�j����~p��UϿ��ܻ{gֵ��&7-��Mnn�?{�-r6�d-MO�W�5�����g�*�ڷK�Љv��&&��1�9l1�q �p�6�Rȥp���`��aQY6�y4i	�Z��/��E���`�K(�A��y���u�ϧSiH"�1��^H�܉}��� �^�A�б�V� 迣W��JSЯB�w������M�.h;"�<�	��S�����&��=J��R�K���k���S�X��=�6��kl>��!@�6l���1�uJO�'3�*��K��Y&Y�9�a�gפ?��4����&�������P���ľ!�ق����ϼ�����u@4gN{�������C[�=�I+�qc��q@;�F�C��ez�����,p���1����FCwL����̻���1�\�凉��?E5IPq��ǡ�tYUi�
�4�r�èc)E��v��M"H��Mz��A*5[�"j�[.���5��6��D���P0I䌭�zm���O6�{�n:����#���?I��	H�dc�6�6ݑ�a�zJJZn�h8cj3O=U#�6<m���:Ȓ�2�`���3��2^W}������h?���f���8��Z����r#'��.O
)�� �ᇷ�U�E�`o4t6��y�"�e�2bJ����n�_ҹ�����(��^�A[���V)֞����6�vJG\�\��r�p
�\*k|�n��㭍�,�.ܶG/�S+(�T�q�I%�}�7�5*5�G��b�m�)�V�2�4hN�^���"�Q.�i�n�6]\�'�,���aYs�Z�o�:��Irs>`��I��xgU�pr��]�=_w�E�K5��=ts��.��N����EGe�F��iY�K����Āv*ʻ���JlO���)������w	�MOFd��~U��.�_A��XpG�e��7Z���d��6~:�����0�۴o�{s�p|#��S	������7�G��R��V�ޞS}�����n�+�n%J��d�J���"(r� 4*oA=��T1J��u���z!ńE���y��T%��^b(	���c���F+���iz1]�LO�5+�]������:]'M,<pT�<���5Er�n"2 ���'N�V����� �:�n�/vQ=V? ~�����b/��ϱ:��b�k��+MhT��2=(����~pf�-6�`�La�^��E4�%HG$G�h'�K��8O\��c���zEY�o�D��#�y�0ط}�݅,7�����W�_��Лc��B���\�o�L��W�zU1�~4Zk�9 ]_F���uU����h�((@6(��LB{?IRL�x?B��S����X*ky\�7�1ɫ��tù�������#���{#�T]e�|vҨ��ۚl�w~��YO6�)˙�B(�CP�;�5[|�_E��u��(�<�U��4Xl�P�m��{���&G⹮X�q�g��0��X]@xq�@B�kJ,l�d�$�x���7��M�~�!Ǿ{��TC�Fe��$ɜ��'Mv�#�?{u��ܖG��7���,3U<�KKv��$!�F� ��TZ�����YЇ��H�ɱ�I��s�K��	�� |,>r�a��g�J�/�bY��?Z�6b���S�^^����hU�d�[����?�z��q���p_�jR�zOe$C	2���;w+׆2����"G�9N���Y �P���s�C1��CjS��}��y�	+X�rOC΁]���� 
o0�Ԝ�i���ω	o��h%C���l�)9 �I�4J�{8�C�0H�t�ࠅ��Ϥnp���[���2�)�Ele�iU�Ç���/#�"�&6ʑz0Q��[wUd�=�Ʌ����,{�K�`����X@��-�VK{�o8f'����_��\'}�=BL�aҰ7��o�u瑘�'���8e3cW����c��s�x�)Q���щP	�5�-T�"���N��2�����V��K�̄̊��S�;_��N�<`p��-|e"��3�M�Mqq��6
,g�Mp7��z�G���W9��̫8\@S��u��2Z�!?^o�����"��i7�$s)�$���Qc�Xz����I=r��;x-5�k�i�
�{؞*6q,�f�R�|K��b�p�{*߆��L�vJ/�	�C�uJN�y���,��A�9;'H��x^*u��I�f�~y�Y�٣��f1�.K��X�B���m�ygE��[�f�,�؍/H���!L�zx~G~��ULwʺk��kL�,�.����tii������w̍�K�Df��G�w2�|�|N�)����'����ʓ�����kEv�\.���xF�ԏD�
���=- ڗ�ގ�@ZP���g<k1.1�&����>�D��� s[��ڟ���+u��jX^��*1�p�aǽ��?���T�r%`���if�Vqġ?�J�}�!���%���j��T�^H�Bț�ƍ"ʁ�sV��Zn�2�/{����]�{�:�;?�	�G`:C�,�+]�Q��.ҧc�������lr�BY�W���owI�G��S2?J(��9<M6QR{T� �E��ظ��{�Ԗh2�
��<�LI��Hѿ�Nh�ű�m�ړ�^���Xr�[`Qb l-�-�m�?H���2k����饘�0�:e��~�ܛO�ۛm�`�SlsN:������اp���Ě3���"�0�L�_�WsOX��1� ����h�@��#E��.�E�oC���M��D��D`�cԾ����#�h`T�4���aPa��ARs/W��#S.��|�i'����j���z�&߮�[��_Ӹ����򾤪�FX�Wן�w�j?��X���������6E���C�j�<��K��̺|D�����k��1�Y
v1�9Yڏ�~�qB�\$�и�E��C�n�L!P+P++�+z�*��῜Ξ�T�/���w�E�f�����
D�NYԐ�g�rQ#X��FTD�s3ufs�1Hr��u�r���*����⵼��D���G28Rȩ[K�=�#�f�$��^u�9(>��7ub�'q���T�����[�l#����vf��9K�lzz���(~^֗z7������U�1/��[+#�/���xM����ə!u���v�C^+��C�2R ӣ�#�:cs$%�/�)��r:y7ɗAG��_��a�(��h�t{̘�J�.u[��W��e�7R�����e�u�� n��]p������v�����ل\ �:�uT�T�چ�L��_��PI=��ΏH�?�0��Nk�@�>��z�&��Jmt�4{���ZPN�5���_���W��^�lb,z�Ţ�l[�S
��iW��y~����c��ڮ����´%�Q�	H��l�6�Ѷ�	�?�z����
D�b�J��UZU��<U�P�[�KS%<�K�#�ҲIv	�V9�ȼԶT��'�p,G���;`��"�][�S?�8�F�!��E�x&w�w߇�n*�xI�2;Gt%o
��d�8f���<�<s{X3q �e};�`�b�[kU��,(g����pq:�!����u�&�b���a��"G��B�8C���koǽ��o��+$�a��F��4�pV�
��6]�� �߆͒��?�n~���>�#��[��2�j��̤�9��~ �!��`�J.5(�.�>�,�0~F�E��I��D�����`=�'~�8Ho7�No���� #{
���8�	��	��HdK)��Z&���!"�BR�v'm�}`���7eaǦ���������q���#`7���g�|90�,��L��a�Yh�)���⣣�`�|�7�N��K�7�{0�F�Zx��j0Tg�]Nq,��q�\�p��,7՗�A���ܒ{2��~Թ�X��`���9x&Kq���C7�|?(��T�a��J�,�W����F�C���"�����hf&�)�^�
FRǕ�nNc���|0��a{����5���r�����,��!z��Y� N������H���H��:6�+��`���}�)��W�dL*鲰��ƛ_�BӶ<v�yL8���v\�������m��T"|�@~�g��%t��yE� ��=�?��n�D>�9�	��q��+ז�������b��%��ݲ^| "����w��C����6d]�[��]JAi�76�H"�h��R���ux' �����%���-���X (T/o�V�>ק[V�?�i�UY��Q`�5�	��ě��^�S��ɪ�<�=>��<1�&�T��9]���y��F�	���s��@�
�� S��_��@y���rJU4�b���߱7�ܢ$9��Q_��HD��㮌��ma"A�1�br=.��)�w)�Tq������P_�b�I�Ë�1#��5�'��f���8�C,C����$y�>�׿E�N���fa�&L���F(f�2\	^����t5`O��pE7	����;{*��Rx��'$ 9�����6��}�O��F��+Q"ya�����_`g�|q��i�1NKn����t�}C��"i��|��A��z�>*�t31i�tO�`m�ip
��Qh�p>����܏M �.���#�*81&䘤�����4F�G�e���CҒ�~T&L�&�4z	�w�pÚ!@k^Q�F�9���P��~a{��v�G��hu��F�t��Rf�H^5�@�ҟ�̎vt���|�0qA��:#9Q��K��<�,Mc���m���3.U�9�NR�i�g��pϚ6���x��u�j�E�7�VK���Z����T�T^]�"K�-�F�[��Y��䟹,&���W���P���ɯ!��`%z}=��n�5ٷ�K��;\�N����=��CGk@�6���47���J^����v��t���nz�`�C�G��cf�8�@@	j�\o`i�ڎ�֭��_� �J4M�1�s��P�lZe+�o��'�iZ��ZkTr:��K��j�{�k�ʛK���������;���>X�b����C+���Hr�h��P.�f�7���')�����Ѳ����c甪�]+ި@5�����>�L�b���P���5�[��ñ�)6��&Is
dN���������������t\�t��٩�_TI,[�o^���O"<`5Rr���聓9��A����<�Nx��7��6��7��/Ⓡ�+��X��y��{�\��t���=`�+��4)�ɜe�c�S��"��(���8�ª�E1+�n��5�aK��P5�C���Q(���`9�lt������/�K�Y���f�M��;k74O�s*�0=M�˽g 訾Ú�|ه��H�K���a�Uu�<��c�4�����c��?�^�u��Fދ���LE�x���č�����'Ν�D�5��>;Z��+�㡠;4�6	�f���V�^Lf���{��79-��| ž��'��Չt���O��&��[a���(N$�����
4ֈk)-���	�R^�zy �_F6��-FЄ�=-�N��KXߤ������b��^��,�R8���Q:$�h� R$�-C���K�[Z����k�L&oW̻��K�U���'�e��C�}}���3�6�C&b���s9 
s~�\kz�� ��wߎ ���JǵQ�	� �b"bl�t���/��1`��?�S�S���1�k���˃"�[�����]�g0U�B�8� r�^S6O�*)~jp����/�#�[6Uq�N5��}��ɇq�p_/�z�P0l8��L�#n9�y�	h�g�L<M�����q7B� �Ə+%�,��<n��B�S�OT�x4�w�H��(b�g�/l�	�&���RL����..�dkn_S��ly���Xp��=�/����^�g�n`a����^*�K�	��N���3P��t��}�,S�܇N��^T;뤟u���C��!�B���6��u�ܜ�s��?��N��uޣ����K�Q����&�E̔h��<rRl���e���2�<�Q�Q"rSp�|3�&ɀ�
�eqn�=�S��K�
�wF�$��`�I��^�����eaFx��*D�7�4�n�L�@�3߂�Gx��$U�P�I?����Ǔ$ʛ�}}�M;~�p5?W���d!��d���AG�
ʷݙ�{��]�Y��:�7/t��M|�=&���{z�����`]de��<��K�j�v���1D�C�Wx9rT���N%+��)w��_:�S������f|�{ޫt��r$X�j�{/ŃA
��o� qV�'wY�o���o���=,�@�*��6(��lL��^�@���Ն��;������|��掚UW�d=-?}$��h�*� ���S	ZA�>�C��������<���BR�St��޽��op"����f�)���B(���6�����0�����I�UM�Mf�҂��J����u�ƫ�+6ߙѰ!bs��{�O�0AKi��^�!�w�ɑd_��[�.���b��8���~�CU@P�kًĳ��o������?I6��Y�]ܵu�9�La8O��G�C�k�=�_�M���C�b�ʂ�c��9���ޠ��.�����Y�S� �� c�X����T�d�{�� �r��=+�g���v��D�k\p�9C��h0���eo6��r��1	,��b���؆>��I~iJJ�Z��C�2�<X����1�W8��~'(q L��4�貽Qճ�Q3yË>�J�J�u~��O�^W}#���(�*��|{Ӹ��Af��d���ˑs5�F�I�x}W�g�,M %9�:R)J��m���S
�ֿXjFj���C�ާێ3O4�-�x��s�ye�00��r�aCq���*��4@��@=�F�?��F^�d�bڛB�7�Im��+�uf'�ʛ�!�˝w���k!,� �)"��5��5x��\T&����ɩ��B{pg� ��Ѓ#+.�����2�[OIp~|U4�3��Ʃ�]�׸�!������L��i�,��ϲ0%�%tY��4i�����;���B��t�l��'Va�Z${�� zn@��*�s��v��	^��lv�q�"�"`:�J����t�6$P�qNx-����"}�>��z�<��:<{�A"3φ�@)/h�i�d�q��5���UM��m3t�F�q�쥃Ν���7���n�&�����C���<#|.�4��B�2�u��r�8~�@�Q#ɳq�͓��?&.:l�>�p��uf _�&`m�n6v8� ��?!�����g&B�S��᥸H��/������-�BnA����_��Y�jo/���`�G�ai"u����׀A��*UUj
3 ���í�si	{h b�.���cwl+��<ĩ5Q$'�C���	��*��_{���4�cR͍=����(�"8�V�ճ>g��,�")�y����.�����2��s�d�3���٥ov!s#��*�g� rM���_���AU�<�5ʍ�u�?��=#�(�^�KVeo���g����o<d&���ܪ��� ;�)$�q!���^�[x�0ko���ӽ�0i��T3�n��/_��2�\>&�&�WV]p�
i��DcԞ���Z��:F������
6�p�8�f��4��z�����C��pW������<����DʶqR��e��(U��E
��3PM8��arp3`s�v�%s=�}����F�;�lq���#n�7^�S� I[W���"M��� ��_��h)�ű���3�Y]-���)Z:�8�?*[�7����7��O�ՊV^z�0��PX�5�������/�zk;n��R�:LM����f�;`�VB8(� � ���U��4*��!�ؾ���`���M�̘���g�zS�?�Ho�r w�"�3-g��񱥆=�8# DR�l˄�VB3U c�:�"�Rge4��,s<�5��1t�Q�9W�,"o�J	r@H+��q�H
<WxH��3���۸礪�T*��?,93i�)/13Mj��r@;}hY�A;O����ͰB�����s�B���C+YYn�W�V>A���f,�X����&��'�����'c0/�\�zެ�*�W�h�Y���r7D]��gh�G��Г �M;�vs��L��fe1R�C?Z���	�"o�ج�ǚq+Z/}t�����ڞ�A��&�3�r����t����`�����|����Gg���~��،���q7�S6��uuZؤ�\Ӵ���a�M>�]�^��С8�r��b�2�܂��9=��)(@�	��Ty�漖j(�v��Zo��:u)��f�Mu�#C�_5M�n.U�fQ.%�l(��y��6�,��:�@�l�>� p�hZlS�����Qw��[�i�<�<mkS�}QyytIy���Շ!�剉L�����.]�:QG�Ub�-e�~ߺ��.�P�Ŝ�#��O(�7���D�ȴ.4��8H�➻��#�mGȰG������0��X�<��J*��`ٳR)&�"�+��H�)t5%��d���\����D��워B�J-���5�@a�6{mW�YV��(
E��~u�yH�JR��|���Ⱦ�k�--�4ho/���u�{f�8c����
��©�NS!������9�����]DQ�P�@ɼx��Q�m���h<����w|����6U��-XIZ�ֈ#�ч^?���t b��k5FA�\]��w����:�Č��S~L�AK0��R�
�al� ��|����ߦ�<@A��ϓ�g\�-֔�W��d��w�2��4}�͍'n��T�c�E:>�q�j}��(��ފ�ż�����3.��[k�Yr@nz�@�rZ����C����M��1�ұ���J����g\}�A<��W0aqй��D��\ I��Q}�>t�^�ukV���|��e��m�6�H.~*㍿�>@�zw��	�=�gXb����ʾ��+yS��O���
�<Tf��(����y�f"�C{o�P��6�o9�x�n��Z�fl�Yת�Y��}�.����b���Q���n�-s]s�o��Ᾰ�Y���X+���o��s�׌��YE4��J�?��X<�6�cv_�$2&��/A	z3C�Y��ʸ-hz���S�#�������z�9Ή����t��W�W&0v;�y�y R���Cƣi^W#�-�Ψ��^�����j��\+�ف�$a��ò�\)iT��2Z�|���j�J8�@��yQ�s-�{B"K5?������X��d��	.y9�(ɣ��#�!εAr����>�(�,��&�)�b�n_�=+AH}E���k���b �g�91|��1xp��ؖT�w�k�h(*�)�*kWO��&Pe��e�DY+�+�ŉ<�a�7����j|�70Y�5��^6����P48��J<�xU|�S������{W-��t��� �N�0�Ome �7~��-Q`�U���G�+��G1 J7!\I�o|���$.hד�R�5X����>�no��ABp��킝ֿ�>�u\��p�V6'HjD����Q�}J���Ǿ]����wr�є���%|���������M��W��?�1��s'��&�o�!\�^�$�wr��9������2����-q�k�M$�Ua�~"e�1y�L7�`�L3I���Gڑ�8��y4ɨ��=P��f�>��Nx�s*���?C�3�a��~:�'�M������Ú��e3��,���T�*�� |�_4�@���0�F
?bY��o/yD�J�dy@������(�Ɏ�ŝ�񫎂�"|�����b3G�t������D˩����)�g��tɺ��P��'��M�[p��'N��͡�sTځA酮�u��vLb�\W3Qp�Z�B�a�,� �֭ID�2���Pb�T���TՇ����u"�,y*�͎�U*�ҝF�˔�1�b��B	��ӯ<����6\���+zT8W��n��˓ R\3�.�^�/m���4�)�ysu�T2;���NT^Xk�����
=s�i�ݗ+���k�w\"y�5�$36�8��:�uW���U�p����xd-�aq|u�h�S�x� ��P�t\�|avD��6����D�X!�"0i�qn���uvVU��s���O.+G�ܐ�� ?Jq�z�#�~C��h��-�0^�l&����V���c����$�;�����ș�8�8�A�䞽�>�gPM�؇�y������x�e>����x�i�(���d�L�8A�L�:6!A��,�<�0��P먶��H��J4?&3��h�B�P��jԦO�~���ջ5�)��+Ub�a�`��60bj^&.���!�����=�%`)�Y/n�ĕ��qn��ҝ{Z��krbE��7�,�L��x��>j��
o��h:�1���+o����鵠�)WH�����09�-F���T�U�_��Z��������RS��43��]���U�^����O�R�������މ2��A�G�@
7��I�zԝ�Z�0��L�n���&(��e�֔�_)e�!���Ḅh�o�f��e,�v�,���� ��0���s�ҏ�k;z�!�̎��RϾ!�Ԕtx���ʬL/��X��R��\���R��}�1�E�������m{�٪�bhK��J�(3��kl���������9{p�,·���!��9C��
+R6���������ǪӴ��P@�p��Kkdj@I���j�L9ۀS5��ZR�P-#���p�����h�$&́*�B����:uW�<��Cyz�>�Sؤ�n�A��G	�Pu�q�R�4�)�fx�5���|=<4ɚ������k�
���(�W=#3�ݗ�1'��J�Ͼ�k����5h1�������t�d�}zCYQ�f(2����l\S�������N�zHh K�<+�7��q俌1����,ι��V��=�!���w]0�Cݘ>^�2$^XE�� ���^�:b1�h�X� KF�{���,j��gO%^�f1�`�� S�.�_Q���g�~[�属��	Q⎁��|B!maI\S�^��&!pd�C�X-I�K��<K�����a(;�L���{��Q�!��#��+�v�;��8�m�{o𦨂��4ƃ�:�����D��OTP�����Ы�|ȟ��������gJ�;h⡭r�q�W@�xrI�n.P�R�Ҽ+D96aY���<����ܳ�sשwa�wtK�q�n�=]���ͭ���Q}��XĒ����wrw��	S�2�4���j��2�0��R��k95�֞�Ws&a�*!����ΰ;6}%�Ћ3�����(�v~6���k:�e�GVr��#�~mL�))�O�,fm��r�9c��R��yaS�ڱ���ku(*'(>pCsa�J�/��lÏ��텵7�f��m���ڗ!k��ڡ%�kz������`���Қ�R���GP6��A��P���ցf��(��-k{Y!T�nO3f|ϻv��M�ɳ�������bN-`�������2	� ���%�[��5�D5���������t���~Ttr����h�!��m���)�p�s�����U�r�g53��=7�1� ݈߳�޾��o��7��e�[��|]�wK��J$zt�� �fϯ�Ʃ��J3�w��%�Z'͠�酪����n�~`ϗ��h@�=ǰ>���Sv:����lDď�$�cȺ�̈`��|l����>����������{��SiD.Q��#���ugU#2�X,*�x����y�:�5o�Jӆ(��?
�1�k`ܕ�~��n���v4U��0����07���Zq��1�2F�ښ�;w��nH�yJ�{F�
��kW��]^O�y��`�X�f��P��.(�*M���*���7_}�$Ȇ�+�~�%<��'�+��!�!����yz.!r�(�{��7'�\�Sja�kI��Em=��'Uƿ���aR�C�ޛxC>�&�J�d���O�,����;�,A�E.���R��f��mI�������M��-!o���jQ����[	c��Z	�X�(����c���	�wt!���ϳ����̓ӭ�Y�&b3�=*���Q�M$FAA=J������ ���N����H��sF����c�T	y�ԯ�����%U����!6��'�|�#u9pE0�K\K�x�\\H�	�%H]��q�p6��uw��^T�U8�Fj�'\�����{�8�j��cXGY�bX�0�m�d�䋑��6 ���XlM
5?y\�:��������;E�d#�5n�s{��.���A8�T%����\�0�Uh�_�p��?�%{�����8�D2(e5v��r�I���8o����l �Y��{�B�(.QH����4ۖ�t�9���<Pߐ�%y������1���)T�'���E������*�����-DXSV�扈�\��Ӻ�����4�2S��	B�5-9�5F���a' ��A)��D��8�]�Ñ�p҅�cY���%Ms�~|�A 5ϳ����pگ�����Z`�%�N��e�۳�d�=Z;�i� �����$PߙH�%�i�����q ����J���V K���}��� �4uQ;Gf����B�
�Cp;S��φ�[X�AU����<��}`�W��D|(��R��9NlY� *1�����Q9��/D��Z���(�d3�%#�
2�[�|�v�1J\PhV_��H�9��l
���g�bh�VZ�����yo��Յm�Wi�ީ�J��K^_d���-�JҚm�J��RG�cDwٰQ/��b>�NR,q�e�o(C���.Zv2�p�O:Ҩ�/�*�ow�7\��HHT�����"1C���2M8��?��P�.â ��1����g��vP{��gC�dCHD��aw��7A�ƨ�rjT$����\{������j�ٲf+�{SΚ��ή�����=�����o��{͸Dn%�E�8�k��:)����r݄�9�_������^=��M�L�!�e������Ǌ2>eQ�)#U���z �Ì��]�ׄ@�e��V��?iR,�{xeG9f�7_tJ��u�׆g=2��BT��$z`��D�*��ɩ�I�� ��9|w���t�G�I�ڐ�d�������H�*�D��Z����ѐnBY;��ze�<,׻�yyR���5H�u2�5zu�qѺ�Y��s�������蜂��Y�D?'���4��>�7����M��q[<�q�9�"�F��a�N%��ݳ�٥�z ��H�w����jbǊ�Q����½�u�J��`��U5ר�vv"sNX���������>X�v@�.�>�׆ml��u��h���9}�q�4��t�������LT�FP$&��u�y�q�MHv9PX	Mf��a����t�-gܽ���
p�����#t%ғH"�����GQ촫\�7�~�'��a���+��A�t�r��:��W�+���$9l�2���*�慁�|�X1Ow2>\������-W�W��S����gZ�w"Xިv6[)�H⩳Z:�B^�6�s#�𥉉:V��r�G�5�?1���sK*0�(�x��ؾ$�x�_y���Y�\ �%ظ���Q��ԗ'9��o���y���qH��|b�h���}9ޕ��yf��K(�"m/��2/���E�=R�]QX��]>�tXcǋϊ��S�{������1��'=g�D�u��ة�=PM&��^���"=s���A^�)�b��o�h����o��+wQt#�x��j�`�<�ڱՄML	n�7	�]8[�d�!J@`�b�Izڟ��j!g���oh,/�ģ�ԥ���ȑ��  �]�@�t�J����f[�zV3W�\JJ����[��ӀYyl�O���uň1U2|wUT��f�����qV����G�zW�͛b���/�z��S�i��"<Me��#0���?���Q��%2�VE��"Z�3�z�J��ț��U��7�g��s��i��f���p�Mʨ'$V6�GM�=O��n�@�w�� Ỷ����?U/ך��y�J�[����oqw^q@)�o���I�T�^q�Է<5�w%]KkD@m,r5*�+f�t����Ж-��jc:P��L|Ę�	!J�+���`˓	 �9�
@<P��^�\�jz��6�E>���6�&m/��N�: 8[�Kq�ʹ��@�Lv;-��D����P�e���oB$�Db����Qj���x8�-��hZ:,͜�6�M�����ʝ�������� ���������t����j���l�J͜��p�9�0� �|���Z`%��j���N#�������b�W�֎�9�A~���;�`���}�a�D���x�Y���0�З�֩�f��pl��rw�|/n��d��J��!GN��#S�����a�֟ɂ�.�9�jr��UHB5H@F��n�帗�ւ�S`*�5�4i Pok��79���E<��H�H`���R^)9R�y]�h�k��v�4V~��7�;[A胀��BW�Y5@��ɑSo���T���󉒒Ǆ�T_�_��yv�����$K�cN?�<���K���ďpȣ�?����@��d��'����-�m��"��J�~������b �x*1�ܦ4�1�Ϥ�C1��mI�ߧ��d�@�I%�H?ՒA�f1k�}Ib�!�3b�ݣ�zJ����؂���r������@�2�٠���k�6�b�v�5���U )8Cc��V?���ҞW���$Oq���c|���v�S�up�����B���Pi>}s����3�K����=��'m�|/�q�n{����WȞ�AX�ї�NQ?G�Z@ڏ$��2%�e���V��:�At��Z��=6�.D]�r��4N�δe�<ϊ��p<4�y�.���1��f����j2*��ҚO_��ɷ�Ww^��~�.&���/�ވZb>Ї�Tc�A�~��߷n[t`ߕ��%�}�����c�,��Z*\�+����&���ME=*n��{�m{�g���*8��A	���i������͓�{0�y�+��ܥv9f2����#x��z	���������!�la��[���dyp^P���k\��{�H�1 "Ύ�U�00zP��)B�i�KP9�����F�眚���S�����,w�6f�3{i��^z]X�Y@��ޮ,S2L�R��W}�)�3|h���ނ%X1ڔ�}=�x�e�$(�4�Q�;2iM;���L����t(aV_�t�d �W�<4���,�������^^a�f����;7�ES	z8]�G�n��H�$��%���ؔ�bE�	���#�%�+�|�5���Y���$���?G��ec3~�d�X�4�ż��hUy���0����r��³)R���]����4(�ͺ�!3^q�1V��	�����\�yjRt��ANHP��xa�� HY3���1��s��ݱ�z[����l��p8��1F.�v�b~I�p����C�Q�]U���:� I8�OH�2�q~:F���J��.�����pӕ���C����5[�/!��ӅI6���3�.��Н����������~>���B��6�Q"�w��k�}@Wv�,3�f�_EB�(��$Ë���:.���W;�IZ.g�ݯh`����r�����u��PJ���� �+Tm����|q�0E��,�����U��1$%��Qb1
��m6� vD��k>P��ц�.�n����e��ЗǞ"^J%��RN���~ё�����̹2�d��d���N��<앐��[@�҄]7�a�i4���˝=\�ԗWDxbj�ը���.�-�#jQ������ń��̣ɱ��au����>"���P,J�U@{�l)���	9Z�$�o�E�%��&1��7��}�Ȱ*�7�!뜈H��ʦ_4h��?/���?��z���B��n-�Fd~��Aha�*Q�_KP8��qnwHI��~���}ڈ^X5���ֱћ35�'�)�[v.Q?�Ml���A���58 �~��d!�ɨބ�P�U��ż�X2+ċ�uf���}@+$�c�Q���� �D�Yԗ���x/+¶�R:Rx�F�t��Ճ�������E�s|���;u��<�:�a�)�)�A�tdR$����`.&OI��y�]��zIuJ�ukES�e�7"����L���4������͢^����-I�=�Q�j��&�:q �
��i���2�"sp����(۸��%�^�H��`eQ�סk��������?�������3�y�����3�ñ7�D��n��RL|�{�О�UL��+�W2C����S��fq�YL��:6'����ܩ��8��|�Rʦ `�F�M��%�f.�D�2)E��+~�]i�h(\G��Lv��Z*��Ҟ�������g��/�L�Մ[�JCKy��]]݃wW	N��<��:�r����:�>��{�)Bo��h�H�e�N�6ɪ鮘Į,?Z�Ƶ���b:�\�a��kBF�����59!���&�U�+j��8D ����%x�ڤ!�y?�΍��� q�~Q��0^0�^�Ɇ%O:"�M�h�������Y�(%i�}��)��B���S'�֖�SK�q���t���,���^8Y��1�Qy�E�&����?&��]�n�ѷ!�7�Q����{s�	���>�z�A�)ǽV��r!��S�k:>����`0c�`��x]��o�'FӕNrIVSDd�3��+�.�c&�6���n}��&���2�`��?=��%�����"��S?�1ǃ�CLFZ�p�S�������;���� ;�m|m=p$��~(��,XS��+<a��Di<�<g��*�r\����'��qPS��.�菒���ա��Bߋ͜��,��aF� �({�]� +uOt��jE����rA]�I{�N�����H]5ߓ0�*o���>]6»�+��e�0�67��Lު�1�j#�T4��GD9n��*����3@p��&�VVҿW��C�o5�{�%�6�yJ�_sku�)�_��\ĉ窠|���7��꺿��S-��Pڨ�߸N�)�ڈK�C�YI�₲�ϧ�=A�=2�5�+wk�O�B�]��Mr(#`��hq%��q�,_?�t
Z���0�t%oI#9�&��q�;(������[#��W��42�C=̦�7��䪎�<�Ĥʂ�tZW�N>�%��b(���C_)�0alL���UO�����O�&Q�)�JD���B��;�t3�K��|�qդ��[|{�
'_��4.=]�B��$���E}D2�-ޯ k��'���~֪�U(|�K��-�C���i�U(��Xؒ�~�L��.2
���z�H��&�OQ+Mu�u�CG?wݑmad��%-�~y=�(�#=�� ��Z�{f�ȹ��[���t(z�-^x��.�CMd��!s~����?��y41��k.�\Dj�2�1DE�w�O�g�3(#�	�9?���3���fG0�b6��tz�=R a��ң`= �֕�ԏ���zw�6�Ǿ�h���D=�����&���(o�>@��a�vݶx��Γ+@8 I�qd�S��O�9#�=\*����Nd<����Q[w#a�S2���
�	إ`G�	��5�b1Lej-�s��͌Уqs����m��F�����J����O;�g�\u[:@A�X��
x�l��""���(���ɨo�x;����8��yJG�#��BD��Mt�Ba��Dn'�b�����a���l��k���	~��ݣ� J�8,��zK�F �9��MI\�Yi�������@w��0S^��Y552ݥ�J� �xfզ1,ld����c&z�<�{b���.�Mv	���윁rF[��½� ŻnVi�$J�s�������.P�{���g��j��3�j�@o������:%tZ)9�I ,�yܭv�hgHX)�	����?Xux�o�Rc��K"܇�h����5�}�$*Zk����T�>l��+ϻFM�[w\B�����!�<��
'�2�:��+^��6�X�`4z"�Σ3G�	�jg @4�lC�㖤łDa�xP+�g}����)��}� ;���w<��h���{wAZ�x�����6���Y�f=H�~�}���.h�K���\�,e��h(��x�[0m�&�6#����.�T�����;���O�)�������
�G�Z(��=l?�}�:c��&m���#M�ZBRx"Zh4�Y?vxUG$�V�_%��ֽ�u�hB�
R���W8���~`"�S2f���H�lǒ��n� <�e�_�P.'(W�f�n�`?�}H�L���T�oh��H�3?=�=�2����J9[q$���)�tm�y#�[SV�����s����NGxuX��������w���V�ԕD48./ʝC_m��^ �t,�F���I��jf${ʕmBXB5�g�J\����x@��w����^h3�t�e��JԄ����R��[:`����bE������/ќ�	]3��?��1=�E@]��u���B����	��l�N���<���""N�CaV�4���[ML>q�T���Fo����@u����1���~l��F����i�oWN�y�"<U���}(�*ZʝWkVD ���3��	������LȻ3�6h�T�b�Ves1�vrjf�x�(�-pq�zA,gD�XV+?�ǔQ��i�������U߀{s��ho'��G�joG�?���3����FM�$\� B��uY��J�"�e�m\��'�~$0-*�ɍz�qvZl0
�-��_܈�!�|�:����A�O'Y�4^��gAn�J�XY�G0&��T����=��ȝ�Ep?��ӊ�R��G� �A�S�\��+LcQA)��uz*�^�*�31Cг|�g���!�I3"�u��/5[�"a�w��1^�&�t��Z}�%.۔Aۤ�����{Պ0N��)���T���[4^G�͖>�}kߢ�r85cI�Nt�ԻB���U@�!�^���0��C��1Bx딀Y���A�}v'��tvnP��|����;����9R4�wl���R�so�RpT$��'P�5'9QE8��PF����ƀ*���(��ڤ[����C�6�)�ũ�P�r����]��W;KhT[�m���m�C�$�?��Q7������	<�'�[���#Wl]�h+�?��Q����_��ccGf�����˔
r?^�}q�䥓TB2xy�&Ȣ`_L���J$��&0�k�A�5��F�Τ<���~ʽԨ���w3���(G����]X&�2
�����i<K�$�,h>���6O���� ;f1��k=Z�;е �q��.=�}wd�&cb����rj���>&�J��~C�NF��W���/��ќn�ҽ�Z�ig��G�B��%���)�gC��
�p`���
�����ҥcE�PVu�#nrK}/br3j�|�z�<�a��PV��K�h��]B�f���&�u�U��X�5o>.aXLg�\�C��9yk&�n	;���4�_'
p=snc���ihDa�/�kѡ��#tA���<.V=�d�HN����|�0�'�A��"oIsٹi��5s@�1�Ds?Q�$�k���P�X�P��4s�.�p���O�D�M0z�3��Q�!�/wB�Gz��28�}���a9�ZB���?�Mh��0�+�U�����9�2iJY�����6J��`������,e�Z1R#��[qnyXh�NY�\1�/��/H,!�G����1l5~$���=��O�i��%D��,�\�V�P�Ś��ipA�$��;Obuu'�,�?	nɑ�=C�N�KV{������9��� ��#�tXs���|��������ͻ�z[����* Z/A8�@%�`�"�O�ر�5�V�U��41��}]BO��H�i�����"��k�;0g�Rr#���nl�\nj$�8+l8��^�]f"1�	��`;-��
����5*�qR��$FF����3���Сz��D�����';�Q�P�̠�"c�0���2��ٳ��G�T��j���*{��� d���Y�T��E|�R�_��6��ڢ]�ݪ/r�~ ����������y��cӖ����^�H��?�A���}��h e-�`��[�\�y�̷ٌo�>]di%Q@��4?���!������`���O(7�`�t}�3B_J/��C�Z\SΤP3�g�qW��?"�-)�q�@��T ������ϳ�v�������u�F������F
=�[IF���L@�q�����p@j�����@�m��\_�~�KcV�醚�����ۮ~E�� X#�׸BP�O�k��d�EݗKǅ�pT7���M�����qk/Ɵ<l|�mM����{ڜ��������{�;zӣ���m���7@��^��\f�ƛ.��3�~n���tm�O$������=�7V�hL-m-i��8r��azT�pұ���3$B����8�s��L'�W�Ls��W�Yꢸ�I{�4N���C})�Ն���vޘ��ãܒ���f-��W$Z���u2�&�ϙ.���408=��`�7mh��|~]�lV�7(1k�Y8��Kc���Ms�U��YGy�曜;T�j}��2�nT�B+��nf�.��]��tK��B��uNS3�U����,�&d�},NBFP��|.�T0�5Zj
�_ %��� 8����ΏS��/�3�M�U��3�������F�R�a�֜=B�M�� R3�i%������Q�O��b@�2Џ}Tc������8��(i�Y�Z	�����ɶ1E���������Uh%�}�7�5���GU���-��}V>)<9��<��a���<Ǵ��L�Yq�����<~J�tqޯ���J�7�y3\񦺔�aJF���{~U8���"��t�G wC�(fiv/:������T�c)yW��0��0+4i�{��%`l����2��J�W+ �AS���~�cب���s�^2*=�hEV�`��쩒�z���`�xk�e���z�vo���Ue����G��Z�����Jr����1m-y7�|����M��kT&1E�l����H��ߧ�;py���g��oF�G��s�WO��b�O��A�h-���Vlk�u2���J[�y�GR.�f I��k�%oxxK?M%�y�l�������/1c�F^�j`��x�����x�Ϡ�s9ɭh˂���h ���M�\�b�-�<��Ƴ>IW~���k�C��P�Gj4BC��B�0x�_j�g�!�<�`��x9K���=�uG8J-�q���*�ly�D����C|���=X�k;''�٫Gތ�,�S�jO��wgRmD�H����+���:��T�����yk��{ )�4��y�>H�1��0��!u�,ɝ�������q�Nj�r�%�9�C]W��nm�l�+Igq�{�n1�WE�b7�D�p�g��E�6���Cv�zz��sr�������ɝ�)Q��C˵��8��$9��$��I�������t��.nď�0%�d�.?�.�!�zR;�ǐ�.@s�f��3���{SfCyȥ�.b,G�*'��\z��$�n@Â���r<#����ڦe޵�ݖ;b �l6b%Rl����'�>GDL�5���'/�({9S�^R�g���Ċ�5��`�#`�n�B
$B ��S�2#�3�t�Dǉ�S���@���G�C�.���1�!�\���/�X��b'��.'^BKb�F��ޟ��Ċk�k��h5k)\�i�ڮ�8���W�g��MP����,�"��{VJ���Z8���r��p?�����=X\Kg�@���DgB�a������Y�����"��KK2�8�N�f�:�m�)�n_P4&�:�Z�ˋ�:� ���i�������-���9�xI�@��~��a��J~V^q�Y6,����n�?h��S�0ͮ�\/��9f'?(����U�$���s�5>�&��52os�Ҭ�?4o)�y�l�x�����
Lt�-�5���).0q�\?�<���l�M�R�@�>�����J��}�H��hw�YH.Y�[��U\��Z��/�Mq0�����<Q6k<O���"�B����ӂ��ma�ͦp(�U����a̍�c��������į�Vty���@���5z�Â��R25�(m�26sq�#fxM�;`й��!ϩ�@2��Y�U��Rv����Jx;�^憫�oޓ�� 妉}�*.���v�<J������,2��ǫ��A ZeX>z�[�����t ���{�M_�>x����8M�l��	x\Uf��J��5P��#�DEߟ*�x�V�jm�0�)�� ����x���'
�jO'7C��h�����F��Xa�PmTb�����2�k��G����S�&�@K�Η^X��r㌻d���o����B�%#��k���!���f���sd����j�,�cP��M�)�g_�+&�9�ҿc"g�����L{�O��k^)�7�/��L�8�W�xS��Ħ�t�`��)�2C�Q�f��48j�h��䡸�*�>�(�u���ߛ/.M��J�RK�aC�Lʧ eJ��v�F�wK�U�(���r��7:��k��Շ���}.�(��6�v3uM��D����!�V0[�"tD6��HXU��~7�m[�?�+ʕ����#(s��.���� �G�cVhu��oܘf��Д� �_P�:>Ŏ���>�cɪ?Z�zo����:b1�.�(?	������&:�y:Z/���	�@ϒ@��e�KF��7�]W���0}�A��&瞼A�I��z&�D@��U�e)+���3$dq�C	���d�{<W`<���EG�Q���(���\�� ��r��y`IF�,Lg�X�0�e-��F̸p;�J"����r#s�+y`�����	 0l��}�"���T��~���Y#����O�χ[���3�Q�5�9ˎ�YNwI=~smJ���lї���6���B����D3����HX�.Ԓ�r����f�br�/��"}�}P���`vtr岶V�p<[�!!�/@&H�TH��X�s�#�.v�D�R&&D������t]5��'�7�E��H��p��;���^���}�w�Ǭp����k��!~Ƴ=~Y9�R�͆��f�7;j��*�j8��'�3M�)`��w�螰��zb=�$ ��O�"�zL��N>�U�w�� pb�-�Id<ۯ:@�ڮ6�7G���&�z� �ZDѦ�!9������]�l@��\:����a�;���Q@��*3�O������g���"+if��D���d�d�<�Cw�ye��ĴhT�?ա�"���ݿk%���|�V�Y��y����bsg����[���ԝ�(O���w�-��tvέ7y����>Ƴg�1t�^A�eq��J�1�.����1�Ɩ�g�\#����H�n��V�#�B#
6@'(���K<�5��%k��
�V��|�c�C�:֩��G���2�,<�[~��XءA�gb��#���}.S#���P��a�2�A��t\V������pO=+YXԡ�9老��O�i��%#�UQ*3���ms��u�b��N!.;]u�9t� ?�2$�#	m�v�ͼ޳Ɩa�����Ysaɲ)'��\p��[���mPaV�(��k.5#�)	Q���.Fj5�h�9+Uv6��Bc=�t����g�)�h ߱�x�m丨��{�h� Ɛ�U�Fs�������u�)�,�f��/��#~����o͒<����O�c���`B��0�%U��*��:_?�1�,�!W�'�!�'0�u|=	rO̤R/�{������ھa��K��/�~�|�OfR�Kh.|�w�ǻwį���1C���=��_�UT��A�T��Ų��/t=j�uk6�����c�����`sBB*����T���Ȝ7���_�)�}�:'�i�pj���"d�ϰ�WV����T�%�ùp�L�-C�G0�������÷d!���x �v��=��W�VЁ�#ܳ=P=ZQtx�.D� DX��	�1Sc��ҟ)��?��`%ws��
����4%y�zA;%}3��]'@0$5+D�Ϋ ��[����q����S�tp֥�x�O�#�ԙ�"#̺Ao�����gĹ���甆܋}����=(d�8?���:;Erf4�lD6)=�4�ZP��h�sJ�j����d\�*L�+:����v�co���AEp�vn
Y�R���%=z��|G�rٓ�-�r.�tQv���c�.e;���#n0�^����*����Z�[}���z8��8�	�kzs��ӊ�8Wc���MsH��ï��4�Ȟ�
�6�,N�Q'ud��j��bڃQ�G�0lY���R��\mY A��b�S�\�-%8�o�`��RR���oBW�x���D�s^K"9n�$����"�hP�������O+u�S�Be��ٙ�B�XV�r=��߇���EҖ���qz����~�y���'�ۄF�Us���Yn %�'l��}��W�U7z$���8�9�(r	NXrG�� �Y���Tq�nGr���9��2�� �=��ˆ��p�^�ra�k|g֭;u�h�+�D�Fx��ˀ���T�� DȸJۈ�ցޅ�MA��i�5m��b�޶ɶ�'�T��ע�a�T�L�o'b˷k���ghN��DQ�=l��&�&���i�g�'gxO�Ίn:�a�j�����[�n7JG�F�ؙ})��dh�&�5�۔�U�G����Y#�ܟ��(�6�r<�s�Q;_��q@ ��v�U��6�9n�"��	 ���:l�����Z��Ja����{8�J(�](�[��Xq'wڋ��8fc��q�R\K�L�O��E�����-�@�^�)��G'8fZ!C��4��簐��j�:?Y���ȈI�Mj��X�OS)y��>j��h�
~��M�q|/�#�<�ʬ�Q��M[�i����Tf;�,�d�,������W�+}9�l^=�o$l�lY��P��q�g8Y[�F R�ؽ������G� �#��R�JL�#��/S��{:��ڐѬ�����"nW���PU7g�8��r�]Q�k�(�[H�=1e��OIx⠆խ~�*�s�۞	0���l!꿳ا� �E���2��Ev�h|�L�W��:TG�RsN�����R�2������;F*hDB�	�0��r�~�4�7�)��[�֚n/�~��>B�J�F"�6� �B[�����;�h��7v��<��'�p��M��e�����MQ�}q��:p1�d�6?I�~�T7W{>���G9j��@)D�׳��!\G��F�D����-aE�oϷH���#��K�>�Z�����.��{��e��5���_/��v��^�ƣ��n�T�c�t�j:�-�C��o7���N6�O�>JD��Y2�1���xh~O-����'M�`%d����W0���a�T�h	��"�-�{����==�q
)/����˴����y9ҜY7DZ�Z9̖'������_GɅ}B �� ,�d�?�9F>�=w�C\�b�N�8'��A"qk�/2+�M\�
H�G�qKn���עPr��B5�"$�8��1i/��>X�ݬ���w-���7��q���2~�ń�üU����@C���ɸ���� ��F�V�^I���}��мt>��Z�:g�U_.�m�^5O.��8�^�LK;rV��+ʎBb#�;{n�᫤ʅ�T�|�m�@CuƳ�V���:K5��8%�!^d�V>���%-��9�S.-D=���`�V?�+���^�Ӭ��ߙ���9�Bى��M�(���-Bv��j\��$� ,�3���!˖��}���.N�rQ�yD
/R�g85R`}��rq�q��  شg�n��e&�6���o��9���a���tp�6 ���э�ş��5ǯ{�i�*�Xs����ݻ��4�A�p8i��榍�T~EYKۊ��d�x�6Vqp��Z�D�e�D���Ps�RU��+���Pޙvd�8Pdh1D;z
�Q��^�p�̥�蟋,A�t Uj��j�MqѪ{%N�I���$M�����9��z�=��u�2`L��i�VD�m�GbJ`8����ӿ�	y�����b��2��O����RZ����)an�@d�y��1��-�Z��xo���߲D���c���㇗���Oe�U5w����ou�Z�;*�ucv|������bJ#��qUޕ�V� M�7E�n�/;_\��1t�3�t���������g�C����W@�V�4���xkf�����6� ��Ԩm5��-����$�͌dE�$��2AJ=:�ED(^���������Ĳ��w,c?�t���*���%�cL��F����7�.u},�'�S������ϱ{n��C7�Bn�� ��n�V�5�\v�yN:o'�-/�Q2g�c'��޳�<�����z3��9�@�$���iP��9�� ��E* �KLad?
(;�g��R���3�t�xqj!򘲕��?C�|6�`hn_B��ز���sޛ��sx�p��=���=��/Ir����9B|t�E�#��ž`�1k5�l{��~�"�q;ɖvs�u�@� ��8٥�d��x��X�l3�W�6�x����wa~�<>mLd��@؁\�qV����22"q���oA�������B�)	0�z7���(А����4S��̪�6�̷�B�+��eJy��>�Q�7���a�r������E��M��uX!K`���]4�7�.TtXR���~��2[��s���7�@+x�	���*�P*�G>i�k��l�8J��f��(�g��~K<��[wP��p$uB���k�L$�<94����d:���X&<��iψ:���#_�����a�:���ߖ���W�n�sŜj�o	c�$��Lܱ|� ���0��xYB��ƲwR�8)@�����(Q���NV�=C��'`C�<�z��u��� �,)'�{�Z�r}	�ω(6����N�*-��l�ϖ���rb�S6�Q��)�,!y���#8��@)Qy� l�����v�w@�q�94<�"F�+m�-j�n�S<V�
�u���)E����^�˙����L��괫��yU���^Z�g�&�J����嫢=�"Z��K�{�}}ɘ�}��DJk��h�#C�&�_#@ji�H;#�܁�!%�>R6t��I�E OJ�|�Ga����ɼ�(q
��j��KČ�8�Ŭa����%z
���bƼ D����gÐX�k���&�˪(+�jy��t�B�j�������
]��NR�̠*�10m��ބ�d���b�s�CxRԤo�;�J� ����:LW��EI�����U��݈}&���A��J.c&q<�K�����w��A��)U�[�?��ֲp"$������lt��X�k^2\9t��kVf�H�kO��4�U�������V��V`E�X6o/����Jņ��g����
�^J�k���c�)��a�I��3�;R(�hf��]>��QZ|��,���a\S�Ӗ=r�"^F%�z��WO���HvH(y��h�Q���~O�t��\�]��#鵰D8.��zcN�M��΍���+H��
#|���Z�I��|��b���꣉�r�SM�@q	k�Vz�$�SȦDa+���HR,��?;��uZ��r�N��Q�K�8�1��qξE�8���p����8�_c�jBO^��:�J����%D���vr�k����"J��P��y��߾Bp~�GR����7�0?�i!,?*P�k���i�$ߎ�ow���X��@�
i���	���a�9)�֘�<����a
Y��湔y�I�l&ԅ��1f����x��!VZ��jְ�Z��}~����p§�L��;�o��ݯ��7�tA
^D�URH�:@��6XVM�S�\r�?<��_��g/���b�z�Zs�J$�4m2v���֝�\/��kS"�h1�ˊX>�f �Ơ�\������#�*%��d�&C?cݗ�s�N5�h[�"��/=W��Kg��@1x��jU�S��V����%�Rt]�^p9��q�o�m/������s��_ڜI��Ʀ^��td'^�l�W����OFYo.t'x��P�q���)�q���-��@!j�4�P�O&9Ka��F�A0��H��f�<K��]�����~�m�J5XE�����>n7T b�3�z2b	�M$�/�2�qU7ǅ��H� .�Dٖd#.]w��E�p����!񟥝&����/����̇t�F�'�e�;������03�x��\�#��By�E4���cn̾Q�jƖ@<����>��#���i�yu��oZ_��*��Ko�8��e�F-u-���7,�F�[���B� T1n�������ٚ�s��d1�Q��4����y�\0��o�<�`%�p��#��r��9-�3Y������\�(�G玮E%�f'����g��R�-3-�y�L� ��,�vE=�*���+t&P�&/����j׻
Z+�[㗒)��,��^��\b]𿷩�^��C��M��_sϱ���#�z4݄!f�G�Fy��-*0
W�T��;�s�/\�>;<ܠO�q��;�G���3�]��h��4�8D�yS�ћ��f�y�Yӵ����AѣT���=v���D�2%�(�OaaX$�n�DVn'�^S^��^��o�G0Q�[��YeiZ�@���oa{�*o��^�����4�=�.犜;#������b��"�/lKd�Rc!H�e��lE����m�:$@Ua�?nc�#^&e��]>Ԙ8���OE����ؒ���#񉽭��]N#"x!��/�g�U8����N9����S���Wn��rek�����fW��vz��"�+c|��O�p���4�x*��Ҧ���Q�M����� ������3����K��*�Oū:]&m<��n)�x[2�+�J�>�����º<>��d�����H!'�P@l$��KB�`��$�(.JI�`2��kz�k;��k O�]�[{�kO����x�GǸ_�URg�HJR��[	��6NA56� �Q¶�GD����V��k�I۬����2�m3K��0�9Rd���f^+'��d�����<����K�"��	�l�.80����W-�����W|�s%gGcxl��Y�uT6 ��tu[OIf+���@R�}0L�h�0JGpO	�"�i���?M��vL�;Y�Z|�w_��`�� >��UA��uyƂ������Q�.#&{���6������B] ��}|�"%�`=A�k��:%xl�Ʉ�w�1i}K@[J��a�+�H��fb���y�H��T�D�GV������L\x.ա����>�>���yE�^�[-��;Ɲ5y��Ԡ@�<I���mŐ-8K?#�ߙ �	#,���JS�.��%�>��2�1�#Ay#jr��i���,�W֪;��xZβ���QՂ��$;���
�'I�����D��
�M:�*`���ɼ�=�o)�#�����~��I�c0l���9�rq��;��ؔS���qjv�h�Pi�.��^����afe�BX�C��t��M��dŽ��nӧ^�g��m����k@�d��S3�Y��"E�H��F�,�t����ٞC��V��u��&V�B�:���&rm
,C�w�3e�Tɣ0d���*�g��P������߳���B�!���6�����l�D����
�<i=?�3��J��V�?�Fh�P����h�g����\���_v'�h���I������3@���Aҫ�ީ����ɢ��f^�v^3�1��;\u��+��Lc�7�|���jĳ�V�_UabxjķlM�w[��	NQ�.�����V��F0G�]ض�+�8�.�H� }��3�'�b{a:�[3Z���s8ʻ@gan���"���B,+��x�ד�^��ܲ@��C�$���ݴ��ƕ�R�������%6Q),�Y��I�<A�zt�+tv���4�4)2ve�Pp��,��M�Y���`p��r�O���x�A`g�/�#+�فH�^��C�̍R+��(�&Pnt�.�W9��}���8�>/*𡫩�A��A�:@E;���<P�񅉉��-�a�d\ky�%đ����8�Q��bn�1[륫�|i�f�Й��B��3+[o])&�̕K�f�`��������<u�$���]e��1(��0���μ�k
��8�����B�&�z�S��7��	�@��÷4�6�s0k���tڒ�?<���_*�f�d�o�9g�VÝH۬�#팗�np)*G<:~ǯ�{B��!�X�`�� Az�@IBfF�2�%Ui����I���ң��&+HC�)>7��)�(��+��_�[�ݕ���&�����H��"�U&]�3aІK9K44y7@� |�B�To/�ز�� �����~Gp�ʏ����O�o��N
H�Ԫ.ĒRI��7�x��*�{��iݢ�����SV.��;���M
%�q��	\��2mUQhh\f��|��̶��Za4�g>	�� .3��"����?L�����	���ߏ
�Ԗ܉`�3Q�'�G%O��pX���U�\n'1�����lW^���1Hl�����}q,��J�׵��擶���&K8��˱����9+����o,6{�X��n�aA‱݈�*t���x���U�p���������i�ӊ��-rS��a��\!���͎|
��yՀ�p��t�����v�eVl�:=�����Sc�AØY��U��k�����݅j��^�$W��`�Gߘ�{�(���
����@��m�*�$�EQը���K�JHh8�yN��t�P�˓�H5<�����9����*[�OF�Aﻦy�#8�R3D�]��t��%�)��Ti�<����ǲS�੊ʑ)�|��k���ٳvd4��޽^�ǀ���ɇ����\臨����4@#�p
�����`c,y��L.��f�h1����t0�&��{%����l�v^^�/$�l��H����a�q��9 �ȧ��c:	�EzP�v)��i�/��nv8{�U7����ݠ�d��v1;�]�f��}K��n��D;}T	z�7���0rPyP�SE��#"�	;8?Ϭ��>��WO��&�CY��U�)�����Dq��v2�H��9OW���lހA��B7"��Ԇs����_��B��tF���3��ۿ���d>10�#�aė.(
�~|i2�0��l�ǀ������_Zm�6�y�}6�׳��R���/�/g�S�1(*Y�S���:�;���0��p'���|��l:1����)���Y��LT���*v�H5`�m�P����`�cѿ�H�x�O�X�r�%7����!�m� 6+�7[ƣ�έX�x�sj
�~�=�Hۮi��G3�������\�RTi�߀��<��:����~?���0��D�q��
{o[�^.N�T�;o9�e뱈���hT�� �����d��	�-QtI&ǡsµC)Q\�[{�ӆD��嫮�P�>��v�=x��D�r W�����On��0nmWƁ���P���s$���������@J,����
_��֔j�uWY�yaŚk���o�2X^��-"+�OIt�|�bx9F��'���sԷ�]��h���O��!�}r���k�t�~V*���{�D��#�������
H�.lbw*�,���I���CL��q��ݐ[����@7Wˍp���_,�sq���a,�v]�\�����î��RzFa���_���O6(�g6�y0�c�QtǱ��3º6:����y�y*7����uR8�+��j���N��5N��Ʊ�����|�&����"L(=��c����w�����:���W���J�j�
f�����g���8m#`9��Ji�ZJ�O�P�}�#{p�̉\A�)F�C}�1��k��d�@M<��_!n�3��a[�~�����Qޫu�%ܖ�J� �$x�E�V>z ���/Җ���@[V+A?G��!$���VF��Y���%q~�;�\�6��G���^��5�CC�CT��J`2��|���޿@bS�(!�}�Y�{$��<��[%�T��!\(k&�	B�����h�a��MN��}n�5�+$���DѾ0K�>$E'< ��;����5�vR�&a��������{��h��<��K�x���0<�5f[�t$\�-l$�
��Հ�C�����6O��5˱M��~�:ɗ�a�b�((X ����p��<�eFz X�H#�	6���μ�����9�#�*_k�-q�;�N�����4��%��DuȽ�>���˦� �d_I��A���Q���VU&�8v2�����Ȋ.�\�Q��]Єh�Lq���m[���OJ���������P��9Aħ��'��	���C��!��Y�\��b���^�]1H!xSEv�������S�W���©�M��d[���R��HcQei1nŗQS�=l�����jjB�j�[�*��{�-7���-���s.�(:��:�=�G�b"#�PK����lB����>bAP 8#S�Ġh��^[͉�=���b����))�K�h	�h�H���
dT�p6>[�,AgZ���b䭘u�L���;�z�mv���g���<[�U�Rp�99�[v�m
���a����(��h�.Ke���`
���V����I1�p�;plr��Ć��]	�@k�F��U[E�I�-3���"~��ZL�a�-�ݳT&�|����3��H��J[\^�,��j�ZL�v�Թ�-�QTDl��H�gb
�N����v�=�~q�h���,x���ߝF��^B��z!ȖhM���]��C?�����q��-qH��f"�`R���~�q���s��6_��<]�}�e��6�)*ψT�:����DoO'�����!ż�Z5�Wr�m����L�Wg��u7�V�t����:�@<j5��ѿ7�3~�� �c���Ӷ
ބ ��g�#�9�S�O�Y.q����';:�O"����^<���l�Zg�͉�m�xCxc1�P�;�W�@��g�sㄝ�Gp�{V��v�bn��������ʷ��_[��e�� �a�Iz_|�����^]�(VT��	ER�M7:vcf�������Ul��V�RHc"����Yr�KO���Q�)@�0�	r`!n���׆&ӄ��Wqd�i�'��P�|�e����_�J��	W���;��uڤ�/7��}U��\q^��r[(l�%=	$ ��̱�.H�wY�a�5�ņSvR��v}�kL���
�~�����׎f�9<aZ>I�xj�Xf�}������i�ɋ���J��#����CŞ��Ks�C&67�N-��Ϋ��8'���ޝ�j�.)��|�@'G�V���B��k���e{�B�	j92/|�̲��W.��?��ӎy�xm�ފ�3d��sU`��v���(��6s&���$�F;Q6��c3Q6�����as��+-���:�wG�*��UW��*U���M������.��^�z�i�Q��=t_^���`�t�FЋ��a��>��+���?�[ƌ4@�����t���sÏ:p'�U%�����6 �5=#t��4�T;Ɖ�4܈�D�:<��U�,t�ņ����z����[;vؕa�ۯ���x�͹$���|l�9t�߾��b��\jx�� �ȇ�=/U�T��EҫM�)2;���0b��]��Q_��*B_h��ߎ�̙�`'ߕ�������窉X��N"3�����;.>�n�!���.1�lk7�\<,�mef��!A��;�)U�C�.�>�=mrM�o���������/�X��������W��K-���h�vq���j:kV:W�E˟\*���X�����Ы@w.,Hh���jR�Y��)�@Gv��C�)��#E2�uL���O �������a}cb��q˚g+~>jw��Up�Ot�σ��%{�Zo�w��6'ѣID��a֙mU�	�P���i�-��9�6Tcjk.BN���1�J��'ޛ�� �y�P�����M�7e�{�5|�]��h�h�)v�R�e�EO1�Ȣ�����f�Mc8��U)��N{Mzs�Bl
�,h�_������(���J)�>!�U�f�zm��ëQ,x���c`p�j�����)���8��A����4xX9$y�f�e ��6�u3���:�B���X-]�Z��!�l���B��xO��StoL�g���Q�ԙrA:�[��*�˲Cl�h�O3a�Yk���mC#���kwjӮ�)�Ζm�cL���@s�r6h�gsdZ@��!�Ks�2���J�ë�]6v�#P�.*o��KL�������P��#aQpQ��g�)a�B+��4��)��a�S�]��K������������
��\I`a cm�*��x��;��2<�c/�p�XL��d�� d�5�'hT��9�9���<w xK��q���s;�4��OP@�\�6=$|�f����*�ԃ0����}�������l����A���S�jf��Jrފ>x\�9zZ)R�ŵ����y�{���QCE�����e�]Z��&���DN$��Nk����wm����[	4Fb�kn��5�گ>���ࢇ2�}�v?S։�ʋ�� ��Đ=>wL�3z�< �Y��>�\�._�E�n5��/��J��Du�8��F����"�0������Ÿ/�gw}�~�7jF���7Z#�� 4c�;D�q,?+��Sp�e
ޭS ���9|tf���3��K'[O�&��1�+sf�iݡ����,T1����}M ��@�&cs�O|�S����)��9*��Ҷ�B3��Ū{H�~�I���O(4_��3�1.�(�r3���k~-V�L�-,=�H��.� ����z\kj��)J�kcӆDK�d/���jh�U9E��1Y��bV���||�k����up���Q�ǿ���`y)��6��M\�J�_ա�"Q+厡�\�*�ӹS���p��8�ur�S�]@.�N�$jx�X�эƳ�ˊ�z�'��z��x^]C9���f#�Zw�A�Z9pƳ3�қ<�,��e%��5x&:ĭ�>����	��gۚ�#���d�������a��K�S`�a<�-h��tSs>N�I�Ց�wK�}�=�(i�)���M�y�Ǫ�r&q�_0���8�8��F\�+���x��H5v��,f*H>ˮ��ʣ6��!P��#�2}1�_��:(��d�M�����#̮� ��!�L�?{q�9���:�D;�* �lOP�9�J�i�:$���1"h�\Q�����=1޸*e�Ѐ��Od5QZT�q*�$�S,{��r^/:����zO��s�gf|������0i��T�&r4^}!�e����!DҔo��I8i��1��	4n\|����`P��c�Ed̄�쿚i��~���LH?`���etx��u��y�ɢ�e"R��KL�Q��q�u��M�&6�k~䄹�Z�Ǵsq�ĳ'�"�������^T���R��&Ja'u;Ӕf�7U;�D��&#�Ȉ��Ei'�Q��!7p���Zؒ<: Q�W'NW0ؓ1s�X�~s�bj�jY��0�>�<��Y�����K�+:��J�G�\����f���4��.8>�].�/�ؽ.h���3h->�ƚߞ��e�0��a�����l
z3pD{c$�2�t�(��tx\����kx��kG�l5J7*ӽ�Ε;tq�f�~�I���R�/���ۨ�Tkp�H���`����V��[��B�:�-q�+e�� �Zɴ>:�Dd�	Q�+�g��c$O�*M���2�RE4��)��1��a�����Y���1V�R�Z̅�׮Q{ֿ ��g���f,D���Jo5c�f�m�=��u�ާ����[N�E�
Г��*�H��!��p崀�45f��a��6�i��`���8���X��3�����`���i�	p7���G|�=�m���4��{Üâx���+�~0�S��6��sE&[qf���D0��-n��/~]8���I���w%-�P!b�qd���N=,�����VY!	�����@��ױ*����$����x&M�!.��dՊ��$��u�	\��_E��'CGL;�	�ygY��73IFs���N���	{N�:��~	����]l�j��r�͚���np���v���z|�������T��V�+�r��*z�R�#^	H�
u�'b�mA�ۀ� �F���T���(�঑x+��`r��@�9��ϗdܕ��&L�U����\Ҧ��ݠ��h�2��y���&��Y��l��	n���zc_M0�Kc�Χ
򮮢Il�*�4�G���qmT�}��#.�W�������;oM#\�Z�	��ܟ�0���k�a�;�fx�;hǑ};� ��v7�Z���ew�������A�R� ��K�َ��������$�eR��40�s�"�,��P˨q�[�D�k��M� ��ͦ�g�~��n�=Щw�t���z8i�r4��u�G5
'_b<�m0�ڈS#��WP�2Ak���e)��N<,ڇ�J�[�Z�}v��!���G�c���m3����,��6�w��(����H�g�bA�v��]���4M�:�\7�wk�j�����w1�a��Տ��ޙsœ~����XUZ���2RJG�z�����R9���tr��:ڗcL� ����otv
&kR��6��]撇v	`��Nr��F���&�c(�$������]W�k0�h��:A�a��ƀ@1��1A�{��B��z!�ޙ��K�7�a���4�M�{B���k�{o��=���T+R$`���T�aX.BFK���@��`�MT�6\s�� �]\v�0�8�_�r�h|X���&��u��T!��'�w9�!���>l!���a~��n�Q�Vf�Z\�V�`m~/eVH}����lrO�}�(�0!:�HJEv���i��iPA�!Y�����}Dt�b��m�zyY��7Tm��8�A���Z���	�~��n���1�R�U�y0���P,�[��{s�<�O�=�}h-iF���8�)�̑������8-U��Ls��Az$�2Xh6sZy��hv�0j�d���|�#�nN1�=n�Z��l�;y(r�̷w��p�0f�i��?��ݮ�	[�;͛���,���CYeT�&��>C��X͡�/7��Mѐ�S���j��1_AT�I�c�=Y0��D���xmd�V'e�5,��W�P�e���RΓ�arX�b�x{��щb�@���`r��i�E%����ڰnj�&�t�%�Ok�W���ʡ��h��\�qK?ݒNX���vs�,pcQX�D�������e�؂׌%�`2DI�$3��e�=�GL�� ������ur�8\e�u �{e�����=w�D^6����o+7Ʉ����r�-[]���q�k=�l�lڷ�G�O��X5�M���E4MD�<+Vd�F����Y6�I���PV�X�� �f�2�v���m��A�~�2's�k��1�M�~L���j%v�$���u}=!*�e0���	3���:'��'��.��a���h�
1|�m�I���X�vp
���-T/����GՌ��=�PPF����ؐdnfC��?)HGZ�Ӟ�|�?*`��6%%����_���/�ɼ�@��N�z��|1�W��Wk�z�0R��E���O�N�ɕJ�֍-��#hҟ�+�D��Rj�7��h���&���t��J��
&:�QG�~C��/�2x�d����V���uB۝K`�d>�칁�Y�ƿgb<H��҆��B����3�{
��C��.<�AYh���C	s�����2 �K�y��Y�RA��L����%�ia�Aީ~(C<H�R��Ï��o�T'��2�N���A(�	�onS3U}��z�q�=�1�0O!��+�3c<a���'{ȁ�$����v����Jj��e��lB�9&�Mɘ��C�S��jݝ�>N�_�(���d���c(��n ��!Q<mڨq�k��Z�.9��3�����%΍`@U!�y�:�}�,�#8Vu���H�KL�[�����l�������`i$ �к�N�<��r��z����H���C!��U�.�T:��C��}�ed�V��5t|�(+��P�pʀ#����,�����y��V/*fq���-�7L��&,>��`$���k �c��ZH�j9}���S�XS��=����a���P�����F�����cx:5�X�2�����
�6ɢ�CfO�m18D���)>�n�<={_�L2���B�fUς�D�Pc��i|$p��b�U�}M�Kބ%b�ae!rm�=x)�R|\����ϯ�;�7s��T'.X#j���@�*C��֮*��S�Z���ڬ����t+f��fخ^�CN\NԺ�Ҵ�
�q� ���G:�zgk>��+�V�]��/t�|X(h�L���m�����#~�E�g�Nd��F�\!5^}<�Uf����e�ܭ���a,Iz�?��������#�$o5�sE�/C;ɽ��F$ؽع#�\G���{����}Z�CZ%�L��1<�N$Sꔐ$$�G*��
����8t�(W�_�>ȵ�	v�p�{*1O������P}k*�a��R���J�UĐh��_a�3leo��ډ��w&Ux�������Ȇ����9�p�0�}|2�V�����Xm�����\��{��{��A
�_�0��������L�:YN�' I�{E�9ð+��+���!��a:7�I��5���>I |~9*��wVر!�D��k��GW�����'�o.�Ѯ
�t�d�;�"
��X����4b�%=�e�w����RO�ć�m�4�Դ�wO��J<���P��ߕ�c��G�Ru� !�_OhU���#̋�н�(���Rk��1)�����LDv�`�_��B�ש����l�jx���!"i&�#��&��"��
��
�W ìx�A��WԖ�nW�J[��jݹ-B{��ю�0�Y����p��ޢ�B��'���`_�9�lp�d���Ӧl����n���{�ν���C4'��,�̰��6�N�U$�~ncĒB�R�pI��(0�0������8��?8��y")�rs�@U�<��0�?��H��be�\#� ����X�u�Ɨ<�em��_�cUSi]��ȟO�nU� L�R0b��ϯu��;�ߺ�i ���<�s�a1���Ϻ���юE���E�A*x���0��@:?Sc-2�#����x�%���'���]]�䅛�=�8L����s�-������?&X\Š��?�hL��Ө/�_�w^���!�S ��nO 1pf��b�&:J�ɾ��껹���V�M30��i�OX����Lqk�Dc�6���P瑢��(�6�u;����׺�1��H=ӲV�pQ�O�ϡ���v��R,�T|�.WV�.̀rj;X���q/8;��\�a�bz�M�+��u�6kB����/ԓ2ˮD�Ф�u��v�
,#�'_����<=2�Q�{��	� jI���R����|�rgz!RM��0�=o��AaFxj�[CvHd~W�3��Q�>>y�w���^e"v��.�1�s���h[���b�A�/�M���p���ӖO$R���s��;�D�����v�iϑI)�X����sŨ�����r8DD1;d䥖�S�|�R�)93�����g� :��:Tj�tb��HR�.+kr����_ةc�j��ƸH���u�^�HGuD�ɋN��]�CoqbN��������{\�G���Yl>!�]<S)����:�q�3g�e^g\�jE&�(u%��tL�� ��]���"#L,�����I^t�_R<Ћ�{w�X놜к�#���R+��\�V�q�"�JGų�R�!�G�faA�0m�q�V�뉜�)ݧ �M�P�➹]���Z��S�!?&S�y��=#b"iVIn8(�	t�d�OŒ�`�L���wQ40���;b^L��#nr�{�_p-;F3"Ԓj���pZ�!,�o0bf:7%\mP���!��@����{�h���Is݋ws�Z��IEno}�Wԯ�����Vq �TDE���vP�����k_��dgep��BMk�| 6}�e~������� �5�h�	�y�g��Z!OB�Y��u���b5Z�	1?q8�C��7�$���� ���=@�l�W7�@�ӓ�b'�P�G�/.7د���Q�ݰ��?N=B�3��_��p��C�RJ��!�L�ˍ�:n��7u8~2zU�g���ǩ� ���J�#���h�XF�`�ޜ�H�Z������K��U�@�(\��`�sKoT�X
��	T�?�6�o���<�};"�x�4�P����_�3�೦����?f���d�8��f �_�wN-���r�6Ac]?�v�}�a,$c�`�%z��֏���(��r�gcZ�7�
UV�(��Op�l+%�2�k�gj�?��sL$� TJ��3_6���qO!�[�H�VY�p#hn�jmSLQ^� �Q ɧ�c_�>&��Ĳ��u����a~ȿ`;�Ѷ�awR\�Ȧ����觢��y(�w���7R ��l�F��n8f���>���p��BT�U��}�h�%l�@�������ȹ��<q��_���Q�'�J"��AKkb�X��p5�e��A�x!�h@m�P^�����;��G�\�Vb�ֈ����[��ӧ��fi_��Χ���|0t���I%� #2� �rpB�
��A6�K��}�e��wQ��%Llͧs#U���Ruj74TN�M�(?�F}���l��pf6D��PŴC�v|f�yF�Y��Pj�9�1�s�R<�{2'uH��l|=��V��]4�<��;�R>~O��ھ9�p`J�<�А+W�����f3 ]�&����2���X���?����o
݉����(k�)�ɹ=�{��x_?�(w��0��^?����R�+�Lq\G�}�[�Wz^�K�%%\J�^ę�rқ�^���i���b���4����/�F����e�uVN�%��h	�{=�8P�	p�6E��a�a�0=7ڗ�D���!2v���TR,e�7\:T"�K9���]f��:��砫�ݿd�D�p����uVJ|�B����w�HQ����Cd!� �B(�"ҳ���21�����ߑ�l�1�"��W����ʪ -�KQ8U���$�>K2}����e�K,R���[��H����	L}�jbU�%�X�|�U���������*�%��q�;�51�q�L�ji�k���C��E��@���3��)����υYq�n�<�o�%��>����a�U���zJ19^��U��SCNTe�?(�����]Z0�6�=��0F?ݣ�.�d�?�X(ހ�� -�9q�V��$����U{�?p#L��Gmp�i�"HŌ��[,:]��x(F[��Ud�嬔�<=�����#�?6��j�B�ۇ(�/ ��+}�3���34��b*bN��AL�~�)�_�����h�T���Jm�����!����_����ǴB��i��w�WR�yB�5���G#��[�M�!QR-nz13c����7wm���#{�Z	q�R/�jC�y���PHC�R�7�t�Fb����G݋�p`���X`(�2(�F�v{�X�{ Dw��'s���y���r�3�*;�RG�ɍW��\����\�3�@Ph��B����r��pA���S���^��,�Т�)9f�?(Z[�>nb9�:�IZ����TmQ;[P��f�Y�����Vq˻��IY�h�s���e3�sF�1B&�.���]zV,�q���'U���@"3c���@��r�G�K�9{�uK��A���eM��ߔ��N���ʲxZ1ZɈ9���Մc���1�S8���q�$�¡�ĢҨW.ヤ�7�(Xlؙ��~_�8Q��@"�h��I�;���u?��K�v����<r2������K�jӋ0�u\�9�*���Ac��R1,R�\,9��# KX��ebN+L6�D��(����9Hf.�T�h�8�>"ҤO�������@�Wf[*���X*���&�G�^��I��� [{�	�I���}S*:�7x>�s�Q���a1Bނۨ�*�+���މ��J�\�E8(�p�J�8��lZ1W�����z�'�#�
��z���yʭ�PVN��c�~���ӟ�	�����)���T|[U�#��èV�I�$��� �����	)����f"E>��s�u�*� )�|�k��)�x��p��븀 ��oz�S�|=H����:u�ƒ?�;�
K8�Y���xq�����E:HV4x<�H����5��b62���c�r��
��o�-��ਈ>e�k��_�к��S=��A�嗔(���O��h�	��$6�k��^*�y��1���@8�,��酏�0�,[�Љ��K +iH�y(���l@x�X,ݫ���b�E���0�F�9�θ���h�`��h��t�-�Z�)�&J�7pۿd�L�K��$�Ȉe�E�j�Ǵ`�*�R���8��U�k��/�B�����Ղ�:�_�L?���w��cʆ�(��2�K[��?g��~x�s�JZ���:l;6�
�1�C�G�j�oG���'n"n-� ѺMf�ƭQ{�#t�'��},$�74���.�����?-al�vFml5_���L�e��}^o�˪����R��i��ܚK�ط�#�R��jV�G����>ym�ߥhn����t/��@pdR�>���[�h䜉H�_kk]���+x� �rEz�Z��B38z���Ǐ���<����2�f�#"���*�'��f��g��UW�b�B'�[Z��
@��wK�����ĩj^�	T��`%��Q��p�>����R:f7�!/&e�,3x�ջ�=<<�xc����ή�!ȕ�mI�Z�vE�^ǰ̬꩝�e���|7~0��G�W�͛K���yjl1� u'-Q�����)��ˇ�:aa�5�m�����S�:���5�uv��j8 dLFPME+Լ ��%��(���U�ҧŧ21��qk�qr�\Q�B��i�b�-�Rt�8���#��?����QH�O��Giq�EA��d�Vh�y��N8�p�d�J{����?�IZ�.���mߐ����|��d�.�%̃u�,�k�����E��y��n0S���a�r�Չ�ge��a�Kw����b�S����Y�����@��͕�59�h��G��N݋����+�9���
�q4[��0x�mU���	*&N��-9�����S6�_��%���ȕ�������1�gx�˔�q�H(�ۉZc����yF��a��O�i}c�(�8"�/4�a��Yq�3ӱ�X� ����E���-{E�A�73����*��j����^�r2�"
.M�qm:L|s
����d�Q����:c��\Ƕ��X�VÙ$��5
'}����vc�����j\�tMKY��w�&�d䞥��,Z�":J�"C����ӷq�*#akލw˕m3S�d��s��34
j��ܱ{Ĝ��n�|�(M#��NB�	%�P�Q�]�xr�kx���"r=[�������V�~"T��/Ѷ|�43B�y����z>��"��Z���/�U��/k\��H��T�A0�z�?�C%#�G��p)DHݞ�5&�� ]FU%��I6��eɷ���2ڢ�_^U�t�۳υC���&)��kgT.�vi����%���r�z[��1�g�0H�� /ϥ+�V���l9"���)�M���I7���0�\\�����_�Ô|Q��L����T��ie��=W �d��p�3U'L�RE��t�����Ⱦ���2փl��P���tn��{"�]���s�r�Ӄt ��g�V$� �TOZ�1h���μ\�Qu;<��uπl�6���n�ӆ:AV6����Ӱ���R�`3����E��id�yݪ��t-�/C	y��7���4k!�`ٕcgw�I�;�٣C*?���,����q)�Svcr-;\G8��F��*��zѧ"sn�U! �졑�Ƣ�=\ɖV�Ӑ�ڗ>��uRfN��":�C�:��)��r�9Ɏ>������?�`R���(߰�M�k#����I%7��o���ڏ,#)>
yE���To�]&K1���G�)d�_��h�!�P�Mm%�ږ��g��9���I���
߇~�5��y�C��i�[O���t,z�J�r ��w����xH^�@���0"�q�->g2�G&@j48;ʍ9�ދ����^��|�6�T=�����]�5}�e�jW� ��(�4W���ڦ���@~��m�PWy[}�O�������Qv-���zKm���ª���/^��7i@+�[ )�؈��/o�^.kh~���{1��̫D]���w��È����xo� �u)���0)j���H)\�����0� 1|@�ʯW[Ͼ��r�n�cz��D����r������.���b7��B2�)9����z"�
/7���N�\;%E%�5)?P���;���~�b��(�L����F.He}��NY�@�	�b6	z��F�c)x7��рi�;�7o�]$��ls�+U�p� ɲ�3W�����B��#��<�iY�p���û�]�6x�$�Un�?,{|��$��fvzc^���Um��.ڧ{G1ӡ���C>�E�C��6!�^u{�V�&9X��P���4F#ŀ�t�.ٺ�Pkuq͖3B����K�˅t�w�/?oH�Ĭ'P���� ڂ�/FJ#���u�KIb�h�3A���(ĝ��1�jo�7��,mV��SF��<9�%��� ,�Ve���D�#T%7��Ӆ�?�J�ē�co{���p�{��=�7��tH_T�,����Cq�9Aurh#r�پO��L�6>��3�U8X��܈X?�j�z����(�JT9��cSʨc��˶��������VbI��%�MW���͢�=���:�W��zL0�Md4OK0�N�ᠿ�_
�N��j?�i�����K�?��(xh2�O.3�꫾JT�]� $��W+�F�?ٌs�/ZLz����d0}8�F<�f9�3��]m�Y�m+�B%�O	���Уؓp���ݓ�}GIc�s��t�wy\��eq-�s��{^��>�>J��lxJ0JrR�8��MO;q���&��=���X��vn����m��7���)�玍�2%�^D3}C�'һ?�Ȕ@��.�Ҡ�i�]z{���Ful���r�i��q'�q[ah?�m��~%���|�gD�O	���f�Sp���!�	�3U��ה��3�ډZ3̆來Z�c\~��uej�`�G�QD"�H΄ǌ����zn��<�[ܖ�W�8~�*����\�Jl�)+�b��J1�>C�9�Im���a�è�$�d�v�]윞�Y�N�Y>x��`1�D~�I�|v�=��8PH���s�ol��q/�WE@�@ٸo�Cn������^��oG["4`>G��$ 8}�)��(�Px��k��S��2�归-�06�+%��w2��ks�E"<hy����F��b�~�4��
�.�p�:+�B�x�?3����8�7I����=!;L��J��!�0I�����q�ECwX��i\yz�����n5�3C:Ȝwu�QR�����X	�½ʅ0�*����t��d�RJ���$�s��W�Za�
�J�'g�q'ܿ�>�	|a�e�:�]��?�`J��"\��O���j����+�Y$�1FJ{�N����E��-�ϵ9&ZO,|vq�bk��δմ��P����H�����ML��a����\G���(���*O�D���W����(���%ڛ{��Y����k Z�"֜E�T��Σ`(x���/���`�ל��x��-;�M��O�E����i���e�},<i>4,��쫣c�����a��8�������<?a�y_іl�w��rK!���'�w����I���Z�z���H�}���})q�떘>fX�Ju���&�[�D��<�zԤ���<����/�`P�y��(�j�z�ֲЇy9�ka���E�����F���4�6by�=��_Z�ޘ��]'S���BRD�..8���[�ξ�Se����]ec%�H��x��t�m����ʺ=D1H����+O��Rab�B�=#����nq��+:������߱C�g0�WI�R�R�Ω�Mf0(C;6V5p��R���	�Ad��=����ȕ[�*�l�y���QK�瑓��� ��O��� ?�T�9E�朠��ef�|�Ϟ�WҌ��N%�P$�GM�#EM>��Ry����)�:PlB��^[}���`�	T�Y�2�[(2$��;,�4����Ļ%�^hҎ��u���PY�K��e�>�'zK����T���ċ�B�)�0��cJ����0��]�z��>�+־֟.���E\\r�����H��Nm�=��p��Y�Aa[e��g�t���B��'�,�|]���~�gM%����LO*]��;�[l��uB|�0U���V�1�����Yvl�H�-zZ+@��S��.��^�O�)�H�i����^���Մk���h�w-m`���>��,-2�9�3;�qE�q��hSF�b�yJ����,�/tp��fBx6-^m|�ζ���a,52����e���jb��$�d��=���|��4\�8~Z�6����e�0�ͨ?���o6�|���h�槠܆����L�WL����x|_���r>E���[(v?��U�F%b���2��;dWk�/	ѐu뚎s��s(�y=�GI_ȼHm'�������а~8�Rq9+��j�aR0��e���"�X�&Z�0��7,��s!oR�g�dx�M%x���al�)QQ�c�~N-��#y��d��mrMO����)��t�5�c�iv��1&�[����zǳ7��b�ɐ!����y��S?� �޸2@J�K�E�hz4�5�h�o��s,E2|K��4��.���If���A�쌔Ÿ��
'A�ᥲI�Q�V��+<��4@ڲZ�,v�;�6���|,F$+;�z?B�q�äs����P̔������n���搡�;�57���,�pA �;YM�:��̡�uI�ɴo��<������
̆�������h��,%�w�|��<-�j�Q%�¾��ζ ���Y������U�+�#����m3<O6���x�K!éV�.�h��[�Ҕ��lK�Ŀ�9���$���(Gr�,�B7S��(驕}�?���3ў��%�C�M�;$���m:'�W�;#Q�8����������I�DIC�ŵ.JQ��N��J��k� Pʚ���!�[j4��ZŃÍWC�_��]i���#TȂ(���Yǟ���r��=�����|�i�3RMm\w˅D�Ց@E��1�6� �=A��R&C���j!�"o@'L�/u�!����}e"zcgWL���J�T�{�'t]8';`b�8�s|�U�j���lm���qk"zQ#r��D�N���x!7�"f3�d�Od�;V��^�!���Vl�8�=N�����瘇��JSe�%�D>c��]5�����QP��MZcu��2@��J�I�HS���J��.���GZY���(����� #%PQ���ZQ�d��R`z�`�)����_*�nu��f�6o+��D0�j�����#SI�Ǟ�t���/g�[cY����欳|ʛ����M�vNT0�t{!���� J��4��nkÝ�-�^d��Ѣ�3~���J]���Ѝ��h�_ɛ��+K�4 �rz��]�Ŷ�+a���Y��*�T�}�I���G�h�4��=(.p�]�&3޴L���CΖZ?��.��`���Dd:U�i4y�����sԨ1~o�l����.Q+�Θ	?t��s�k��s�=산�$�Yd�=P����;���٦�V�;L��w`����v��y�v�0ߪRgV�x@�)׳���+� y�b�������?����50n�Y}�xv.��[ ԡ�~yk�C��YR�^s��J��@��۲z6�9��@����` ����{���LM�x��a^�t�7�U�����,��;�Y��ْԍ_��t3w~�����mX|K@
SD�\�M7N�"�؀w�����RF��[���
�Q���|�v	4R3�@�z�,{�3
~t@�Bژ��o��M`R���U��������E�m5�S0Os��y1�]L�u���j�}Y��ES��/{�w��(�9�[��I>�C.�\���6lE�H��o�/T��c���V�^�X�:�d@QZ�u��e8T�G�d��AqP벱/�(eh��F%���P����c6r*9]\�X��6!�3NT�6�l��;)�7)�~�l��E�(�cUf���fW7������ZHK������P��f�KGz�����O/�9��^e�mW޴S�T}x������*�7�Q��Ⱦq�5���][��Ƣ��jƁ��+���Z�?��@�̚������s-����BU�Vsq\�Q���1����"�"2��K�$8�)�Nb$|��Ĩ%���V{��Ri#S�������9�y�p���r�b>��dyҞYaA�� :�%$��L�*1����v��E	<�������I2:I�]�粤^�4A	e� ^l��Lc��:{4n�0��D�|旂��y�;l��h�	���t��TNʺ|%���3��V�����<�7ktem�q�I�%Q�ܟ~Oz����jQY������߰,�lO	�"�+�
�f{��E%���+� �&��	ǹmx1M��!b�-A�׭��n��������ds��m��,]��/�i��6��W�����A��Q����VN
Yp$w�g�߷s�K��H��`[�k� b�λ��-�E���ۙ���W�+���~��]���7g��?A�u�f�'mV��Ö��UoD/����Iۇ x{)�J1�'ݵ��g$�:�z��H�4�S@T������.�.�t��l�&Pa���4���T�wH���W9�L�D��������5:��E�W<G©�n���;$����J3[㤖��m!�̃3�����C��%�qL�ۉ���{���	c�*����4�(�	���1;�E@�)P��o�i�x$�L� +�K�Cd{�&�S3h��6P��]r1�?�ƶ.�f��Qt���w>����dm�8}�i"��֐&,��4��H�5^!&�e�o&	�gB���.�"����J$�"�PF{� .Z|������Z�^���4,fؑ\��N\	^��6�-{A��U�V%h.\,Ͷ����N����偖�ǫ��Lل]k';:��7�1�eJv#�����ƫ��F�Kpr�FO-��ز�	bz/��G�F��>ᥘ�J�Fd�E��MS7�o�:&�?�2E� �C�d�+�񚑒�7�4>&f����v6��7����������ML뀰����w�tH[�!���<,df��j+��d�`�����އ������3鐺w�:�O����'�,/OzY�P�o�eT0y#��n��vQ�C-k)�~1�fkY�.2��$n��3�F�7���+�Zz�+C���6���F��qe�u����h�dSA���j�|��{;bF��!Hm�ra���q���r��ŭ�+��
hr�?T�$�	6��i���z!�%k'�#�y��I~��B�&Ǒ�^��)ر�
�U^!���a\ʤ�ַ�͡1q+��m!�4v"P$��̀t@eg���.�clRأ)ĺ��^4�c����y�h�kKP��0,���*��Va�*��dMsF�	^�2	YBd��UDd��ov���)�=�N�u����ƭ^��kF����2�w0��C7@k�t����d�(Ef�eu5���`�xzd[p�?�]��t3f��4�𩵫p[�)y����?
�G�dA�r��x~@���AxmL���E��@Q5�'�V�VW�T%
�����:t���������h$qAN� zʬJ�B#t���j�]��6=���5���ypM ���\�r����thQ�q:>�ƗR��
]��Y�?y_2E"}��0TRƚ��P�3t��|�`�W=g�F����3Uڐ���sǐ���Yn�<YB�˸�'Aދyp.�x�<�J� y2�Tcp�0c�Z�Vr%
"��ܛ|�I����>�4:�~��v(XH�Vl�j�i�vf�Lv�A�8❘ʀ
�]#YE��/�1�hٺ���)�W6|=�8&w�-�a��ܥ|�L�ًeP�ό�nh��kv�mWɩ@��=Z�;��}�����f��Ğ��cu�d+�67I"���=b���zw�[J2����LIq��*�i�6��>�����_<�4wºyD�0r��~	��j���ƈ��dY����Z3�|�WL6@4:���@�A008�s�����߷�VA�o�����a�͸����H%�s�x��1(�b.�|&�AM-����V�_�w�	�nU�� E�gC��,ӂ�����E� �|�"[�Mk�&Kvԃ�1�;;��֪ 20C m��=�}���p�����H�z��D/�G��e��,�;���Tp/u�����LѰXFG߅-j�7� 
�J����$�͝�W����ݳ}&���#D�Aa�}��`�Zj�|��p>�9��IY[�1p��b�"�,��F��?AM��}f������~�«�ב�S/pR�&}fdz��ZNU#�Ʀ}��k����E�E՞��'��;��������JP!��)b�F6%��E,�N��Q:l��C��)�T�AHT���hO�ȮKn!�"t�x���c���mM8o�,[���H�y����x�D+����Z��~��f��S����Ò|:>�<���pNe0�"�n���l԰<b�2�x�[?��(�#�t"Ѡ_ɟ�JOsT6i�����fw�3��?�D`
�9�>tN�\1�NG�����
$��eHþ.l�H�w��+iP�s�� ´�eH�T���b����Ɯ��RVF��-*5a����ڣ\8@�N��Ϸؠ��qȱ�<Ǎ̞߮H�v�4��<��Q�1�P��4��Ǫ��c�Tݖ��Ba�=�Oe3@����H��"،�=��m��wj��^�rON�"��PG�{���[~�'2��L���h��@�G������Z�=d�L�n�S��:�`вB)�	����-_)-����iv��:�������2Hw^��^�o�{��țg'�g>�^��-l�iq�#
+cM��ڔ�iVQж�=�d�	ξ*��J��=���V�|rdz�����wL�V������Я6�u�q91��F	�Z�AP�ǽ�z��E�C�ԇ�9��xh�������d9Į^H���Že���)���/@�g��� Y�{]�C�����t�G���W�7+��z��#�5�,��ndݿ~m��Ĕ>=�KH}�y���H�����|��Vr�ߧ�n�Y�e�v7����cE�V\�ւ��O������� ���942�����M��M�@���F����aȥQ~[n������t��O��"=��Sl�L����a�Ԃ-.~te���ZQqe[���Lb9��-�h���:y�DU���}���B�-��,�L���W@I	��q�_�O�~.��S���?���:��� \M8��`��z�Y�4U�H
�h�;��#v��e�W���\�vͣ�m����b��N�*���`�/ؠ�}�M7҇ki�s�o����&W��C{��<_V�0&��bV���ՃM[;��b��|?J
��7���}}k�t��z��8E���v��+șL� �g�3�"rj'k�� ,#
����%�c�r��҆�Cw�m�����E\F�<-��Z��Ū��',W��Σ;��*��
�����2�V���7\�q�*|����~��,����z%�*jJ�)u '>����"���p[�@����4d���y�z�}h0<�(�V�;\?ORy<P.`��1������YaP>"H��?����ok8������$�2�?E���k����Y������~�&!r���oW�NVૌM�K�HV
6�0�$�7Po:�f��3�]#����Su��fd���nP��5Z6��<���`Ox����_ތ��B���eq�{L���^�ۨ�zCA�,�5wy�V�ՄK��w�JoQ^ECriu9��z{�a�5S���h<m���h�� )��H:�<=Y^�D�0jt���k3�.!n`�tT�M�Ќwf(�����I�)�(*��s+HN#�b{�x���R×G��WIc�N�0���'@��U���˕��fk\���C	��󈡖pG��Ե2 [��x\0H}+e+qG/�͜�2�m�=Q��ɇR�pDK0��馀]�W'F�_�c�"`��|yQ�ϧ%t���m��D��:��͔��6ѳ����Z�_�v���P|��0T�ߟ ��tS���w����?Qlo�����Ԋ����F��ެ�P�������%ۺ��7�ǛQ�|l�r	<\/Y���pK���0H�VL��& %tg9H���͖OH��LH������#�	�8��h;9��a�oC�[�ݧ��3(l�vG��������=�/�5�S҂���{�$fH��0�%�UO�T��l�Q���h��hf�,{�����.�M����;�o�B|���N8��V��Z+E �B������J��Q�BUIrl�^W�����Ӆ���`���S�q�t|��ܜi���y��bI���Ujl����^./�:k�ki���G �{}/�#��������"���K��Dzg�����D?h�ծ0�U�q�:T��J�K��Y�a�|Y-2	z���?ҝ ������u�����ټe�8y���^�j2R��abQ`�c��W�ۀ)l�G%30���`��<�ٹ�3p���R�Szm̃�����V����J}�(���A�C�7�>W�t]L���,��2�������G}��ie�꿐J�f�ۡ`k�W*�ַ��^��^ؚ:zD�BA�yځë�G{��I/!���&xVp�1��i�� �b��F��A�x񈴭���&_@H ޫ3@n9@��]�4��*Ͽ{f��9��@�"ߓ�D�4)�����s�H�$����4�>��\ab���P)�c��CaI wu]MuB��� �BI9��6]�xC�m�Po�j_����\���s�U������� t�q���)ic#L�Îs�LMX��k]��r���3�ª�FW�K~#C"����c�b�u%|1��	-4o ^�a���%�O��ߵ�# E�j��Ŀ����{����7d[�:�h��{`4� ,X�щ�ѕ��jVپ��ta�ߍ <B@��'�?y�����¢G��T�UX��M(�u�Q�PvL�K���	��p�ΫX}�T~��F��k���a�{Ǻ ��8Z� �K �����X\�����u�s:�7u����s�\��P��甧�R�0a,W��T�;-�Z���^��>�ݨtY��(��ν��,J���`&�x���IG�+�N�tRآu��
�g�(��Q��Sb o�B��H���}k�^w�볆�R��W��c���$���T��t9��K�!��]�� gM���I�Ud^J���K�%��S��DC�d<�ܒ7G�vL�N������C�e��I�.��o2*v�"��f��r�W;IW�H����GI��s^��?��l/p�	��GR�0�uDg���J6���X�I�!����w�o������KV~߻#�>�/�^���_r�s�ƍ�;HǕ�%"�X��`���W���H?�5N�y��*�K��n��0�1�yi#�O����TK�jQb�=#�%��o!埢zo�~x�0WÆʠ�;�O�>�I�9� &��,���������+�2~IB�хD(��7��?�-�����1���!�J����X����p�8\����˴s:��e����u:_�]���*�4(+L��j9c�0�O�v߿n^��E1�q61.<��b�Z7MB��|v��몺�}�O��I��$K�ʈ�U1�~u�caỉ��e�铢�m��]�aI���'.^�DY�4(�
�:��Ѷ_0��s?� g��:)�r��v�&w�o��� ѭG6�E}��^$Z���U�><OҼ˾]�6�Z1���,)�y�>�̎�}�;[(��ސ�>D?���U�v�;��������ue�W���1�2�
�8��)��V�3�,������ԋh���7�i��d!�lY\��-ؽ5�d���͉��ͳ�38F����!�XQ	�b���Z�e�]���M�Y5��cfXA@�()F�ku�(���U�{��@�>
�1)��G��'pq��\�����.����$�j*�ƸČ��f�e��E���.<�ʯ��0��Kݎ�mcl�~��c>p������Q̷�����6��U��6��u��5}tX-F�	y�O�QdѢz�ɽQ���8*�y5s2C�!U��iO���M<������N+ycco*䟧Ǐ޻
�����p����+{�H��$�V��0�%'Dwٚ�R��/�n�=�Cj��d�(��O��y����v��#��������rN�F0�K���@$,�� �![��%g�Ii���'|AK�K���|Q!~���W�EI�<�r�Q�[�=h�����L���"�S�{�O��;xz�3�翬�/>\�����oa�X����0���ӥ#��N�"#Zb��RU�c ��x-��k��эo�קsOfD��8č�6&��B���8��!����͏\�5
�.�ِ"a�>���r�����y��O	 [����y��@3t�ǅ" ��}�ux! _�7�m�nM���-��~�6 @�6�4���|6���������KJ}����TLo�K�,#7B�����:�x��S^W0Ii�@�H
�[	糧u��� Ҙ�,�y�c�	�V�7(��6_v���T����|2��MҤ��b肴�߄�Nb�Q���Έ�k`�e�'4I,t�%-p�U�*eD���6Կ&��j�;��q��Kv���BN��}�E��G\@.e�ky��&�1�U��c*C�*�I��_���v�'�MX�5@<��E�k��%�C��\0�8�3T��P��8�5Oh��uQ�(�z/
"`�o'��1 x@>���g�Е��3���|ɐҖ�\��i�Pţ�������[��9Re[q"�#</;�u��j����"q��?O.��x�IP�=�|[���i���������JIWj�c}D���#�i'��!� ������S	��c�g6�PF����Դ6B�m?'�B}�Z
Ab_�r�ξ���Q@D��$Q�g���ʙӺ���q�Pau}�J��w�4�ɳ>�0i��.1� ��69
ٿ�eG�KU��
�*o
�o��㵞RH�!�v����<K�U�|M��
|�;�DIAd�zg�l���"F���g0��=
s1^wY�X���&&EC�ȁGtK��xms3��??_���$�_� �db���Cm���=b��?SU�G�a"�,���\�e�(k��tVˎ�5H}ץ�A���?��.�5b��O�r*d)վ�N*c���;ugD���"zC)%P� K#��{0:�i�M��Y��	��o��V�s^�PW�w�ط'�n�;�Nx"�9bku�S���v�s�g]�P���4J��k�ڻ�E�V�~�):}葸-��2�3J�F}�2�����phbn�k=$����ڌ���.<'�q������VؘǱ�WC�!� ����������Uɓ��Z�F�y�;��[I5KA���i�7��)�����a�܃��[]�К�)7]T\��b	��m�'����Q`?��L��5��h��"T꟦�Y��fB�ٮP��qj.��'E�&V���.u���T+���=��]#^�����1����X>2��'� �궆���5��FF��R���6�'N_�	�&g*�*�I���3^�_�MF0���&U�1V�D��TJ��!9��0��`�=���u4k%ez��x�~m�g���Z?K_-.u�J[�k��`���N����Cr� 4f
��<w���U��)dϪ ��!!�\?K����`1�+��c=K��p�eF��M��B�M �H�6��GS��j�>]9��*���lhs����v�G�ٺ\�~_�߲H"u��l� .��
�WKA��Ks?E�c���V/	���n�8�~;�[��#����0&4�g~~�u�����?ԩ�����Tf�m�"IV���`6�����{��-�h����"���4�u�1C��s�.�h��ݫAB �a�����i@@�����R	ԄW�q�r��N���V�J�%~+���𶸮;�Mɡ��R��+)q�voʈ5�A��$�-�ϔ�Q͊E@�I�Ɋ���ka�'ϛz�����RH%Bt�	ڟ�}P���ob���i� 
_��Q�U0G�K���sj�u�X@��S�#M�BH��Z�[-��3Xn]��>��N���bb�Hd��-1<��I!�,��JKLTX�PZ��!���s5 3z0"2*�� �#�ͱ+��-;�1�MlJ�
���g^(��k�
�����Oef���
�]ń_��}Di��~@HLb���I�kC맀��d��Uv�#	Rm_3����һLʖ���� ��\��NO��z�Ɖ�W%��n���~�{�s쳭d���W��\"�9�SmNz8�	`���2��^��c��Cʌ+�v����6ic/o:U���;B�^Gʥ���f��ꍍӵ$����l�f���βͰ�u)?]c�馪�{~X���8�-�*w:�)�t=�<��k}���ק�E�3gh�Si���6O� ���jr��H����@ G��Hʚ{�eB/��%�
��Q^��mea�p�e��'ge$^�|��l�[���<6B���p����-���MDZ�g��CmsKF��el�k��wπ|
W`e��}�h��[� �~�����N�q����\��-TCm�(�I�B����-!��P�ȁ7��u+>�f}2h�iВn�u���_��})&�54��;꜃H�@���K1�RBn_��� �X0�K�����}��կn���H�܋[��c�p���^n�Bq��h���B)���^b�c_���+�q*��t��tWKe��C�p��!HB4A�5=�\q��p
�@�V���c6�3X@D|����\U7���� �J���Aٮ������=�;�O�;H�kXaO�@��s��i&��s/�V��rQ8o��FMc�x�9�kSfK���M�xVw��!�¿�ɅGԈ0-=`'!�U�fh.���ǽ�����Pz+��~�Q?���݆��� ��h�Q!cX��0�Q�~�l����6[l���(��Ž��2<-S�M�=bhFQ�D�1>G�uu^��_{���K�3۩i'����
S�WP/��B����T`��㉬�m2�I	Z��S;���n�Fbe]Kc[��;(�hC<SR�\E��(���/�>�}�`��:I�K�ۚ� u%�ƴ�J?�4�{��Wlǃ]�t7�����GC�APf�kg>�_N1��[Ed�=���2�����^TW��2�o��f/�waZ��]O���������L���H�=�)p%A����7�5�k>Y?�-��*���4�S�B@��n�9uw#b>c�#�H��H��Tw�n����.��8�ʓ{s+��	)=id�pP+	�9����׶2�YLԿb؉��8`�g�;�u�ywMm�mF�x�"��\�	R-G>H����b��	��^��|�,B^��>������z�tD���\�R�܄j�s������qX�9�
D�,.e�-�Y.tyά$�<M�+�}���X_>�׻6����R�;�gҚ�g��z1%;bv♻]�z�f/��T�^�P��8V)�)����!�J�F�����۩�~�_.U���fw}�"�:�q%f��'����aV�K��
��������x�'�ހ��������"�pS���:�A �V�cNZG+���ALg��%UrbZ��8@�!�h��L
yx��S9���M@QH]I�0�*"�]��ʻ�ֱ���	>z��'>�i�+S0��N�2�X�3�]�p���3j��T��1�_nN����e��ܐ�H��h�3��#��ۇFO����܀�n���c�AT�_��ԃa|F9��k{���uAJ��y^���qu�l�{6�{��dH8��Bv@\�C_�T,҈�vz�C*�S����}O]i��0@�w�.��V�?��p�P���܎m�K�'�vĊu�x$�|.V�w]g���WV~����53�;��vB��-���*�]����7���p1��E���6��F�P�����N�L���DY/��7�Sʤ<ʟ��w�AM)`D�oR�~L�4�]�H�|���מO��98�3��wQBPx��������(
���WM\�$��/3W3q
��Sw�'�Uj�?#_؆@䘀�bI��j�H�X�����[(~�hu�h@�RЃ1o�ٗ�������玳��_�]i�U���=^�v"tzV^�Ql�∰�y����ܕ�r����N �f3��vs��cQ��EBRda�̣d�ە�q�X�p�dF�I��>H����/~�2�q��U7�0��������>�������r�ip��Pf��o��6s|�J4�R����5�Ŕ��� g�	���p͵�Ci�g4<Ȕ�a�O��z=@1+gilly����ɜ��(S�,,oP���&�q��M�7���	$���¢�i�5�
6��T�<����\�����AI�$����}��Mc�H���ғ5V�49X�E��t���?o�0<�d^�i�N��4Q�O�n�
���{��e'h:�!�����^-�:��b��m����q� �� +�s�O��!�����\x�oq��|.ݣ����W](E)����ͬ�ĀQ��)[֘Ao����CAJ�@�ʔ�:іv�����(m6S��5_M�+ڻ���!������C�B�YP�����:9b�˷��z��8?t�'g�t�%�9n��vi0�`N�����֕�N�ak����/�n?ͿLw���5Rx��d��. H%�QO�+�3�ubx�Y#���XZL�$�M�i�!d�<^ౣ��}�`�i����X�;=e���K��Vn�J2 m�bP�K��Й����
"�kD�B^0=L���;�otk��i�J�}1�|!�z�NRtE&&*5ߒ��rs���Q)/7éS�!�w�'�G��J���]������=4AL�WV\z�v6��������O���S��Yʃ��8^!�j�{�xW�Q�X��1ay�M��YŒ���bb?tF�}Ua�z�?�.U��;�h�$�]�_(��~<7���zw��D�B�ኻkzpM��
�d�����L���B�k�O~��9�짾S|���L�du� #^�xPX��j$�G�6�{Ԩ��o3�� ���D�	��j����\����Yl��7�$7;&2��JK�LD�?�OxAS+%5���B)�;��;�B���M�~�w,�������5(�h��?/V�W�nX�����\֜Eݬ��������̓cC��NcH:�[�����ۊk�}".-�'�,�܈L(?Z��[�׿�}�;{Ÿk�S�5���qNsq��,�_��h.pչ)��M����I�6(k3j���).+�������3#�PPt�.��tô��!�29��	������My��}��'�Y��g;�Fh���X��S�`� =�a$>�Ϛ&#�fu��ʄ,���h�����{�� Ě��>��d�5�b�V���fg�0[��[��b̷�W�mL\ͳ������.��[����E��$9:�$�����N�L�ɀXu�M�{{~~���f�x]d��bSzupRk��ؿˣ仹���g���Mt"�$�Ć�ӦY���X��|ߌ�U�UN�z����i	�6j3Ph�������}*��y5����X�D�R,w���3�P9�*�ۓ$��~DV���Zs�CFN�Y9:�o����Z >&|��{լ/n����ߛ*\�� 3�,.R�j"�	�?�[
IP0��(^d]��:3s�d��L�ŧ���I��é{�T<�eI�N�]ӵ����tf ���'�h]�S%�m���Zl�)CGq��\I�Ǐ�Bt�3X�N�T�h��H� ���ud˂�-�B���&�� 
���TN}�	Z���I��]ol������T� #!H�[��������y�XV��{!�t�-��{��]�{ZR�Dƍx�>�
�pmR��d9?����x��4)Í&���Oq������;��[X����'����3�`�Ʒ�*�9�^cT�����*��"�-�!��Bt����E&���Y��8L#�����y�X5����*��f�Y�k��E��T�%���ڪ[ee�<f˸�z���n�E��P%tw����mK�s�S@!��w��r�q2�������d2��k�c�؛��E����j#�t�9k�afˠ�eŔ.����X*v�����?eJgjcP-ZT�P����t�ycEC�/���c9U0v��隡�5�%��3���*T�P(������$��[���u�)i�d|���_��.��ߢL���]��}�>��NY1J�%�G)� ɹ-9�>��x�ޗ�a���B'�u�w�{�vǪ�',i�%f�*��4�g&#mP��9%Ǆ�|��R��Հ���"yv���fi?+�u�������4�Dx���|��eU�yJ�*Ҕ�LC)���%<��+�y�v$�}0��@˯'=N!�g�Tϳ�©w�:=�u��H !�K��4g����?S�B<D��2!�Ɓ�	�ZϰoLϛ��0o�z��M�⭾�'�lt�xb�̩�G�~f6�Rݼ����f�ig*	12�Puƪ,1�D��(z"�@��^~8H��y�e�iCKY����B����Ѐ���l��R�Wy-�܋5�W��SCWn����&���8�%��]��x���i�5>Õ-�?�xy[��z�_J/َu��rM�#ZR����nnr5?k�q��hx>��P��;�ֵ����+�[KΌrD��d��4[7-��:�'�
�=;�Wh]J��`>ZВ�N��M�Z*͵=� ne��`��P�����q��d�gr ����a����>m��z�&�.��9q��z�v��e�_kY�ic�s�T	z"��=�3��������l��gyp�|n��ς���IG�z`m��c)joƁ�8=��]�al����ÿ6��������l�\�W���&q]!f�H�cO���Έ胳���<�5�RX��|�Yʽ+�6}I���cD�d���Hm	��8�%�0��TCj�&��k���h�	��g���G�q�LL�*� n<@┇~�,Jw���83)gm��z�e�+���db4�Cu��{�wW���Y�&�hPq����V���r?_*��=P&M���ISM�Xk C�i	% �]��Ş|z�2�1A�%��K����}ݺvo�B�h��K%\$�Ԛ�H"a�ϰ0{v|��ℤ@ �M{�N K�^�<�$��Q����M�:y������]z��v1�F�`@5�<ΗFo�^6�R�-޿��욢�K1Mv2q�uO��a�!c[��Kف�΀xF���W^K~�2-U�)��ӗɰ�����r	���}��]�忱n���5�J����GH�6]�{��%�i�t ��R!O���i�Hg�g衮����6�l�m�X	��W��J�)ጪ��}ڣ5'CL�S��y�������JT�%����^!���I� �����Yq�7q�Y�<�`3��e;����(�Zl]K�LL�`6f^�!7o�5�l���A�����ܫ�7d�(�t%�-� V�# g���I��c"�)�P� 	#�T��ӄ�����β,{�*	�d���h���L��.�}���J ��J��̞�s�|џ�?{a�'�jǤ1��:6%�������/�kv�"]���d���+���b�A�����"G.1;x��E&��ǅ5v���~�_����T�:g,c��� yȈ<N��s�1�~Ψ��z��\�_�
�Y�}��z���Am_<��<����Qr�@d�#�Ћ��H�R��b����L����%�4���/�4��0��l��"S�rN�[8�-l����V�CѲ��T�'�I"S�׺4��0�;�t�Lb���s�nx:�m��|(+��5���J�g����*s�&�*�����S����4�kq�}�w���ZLmS�]T�[Z�h��/��g�ƾ,���qe(8��"
�	.�l����e��쀘��\դW�����Κ���oK�U@kM�����%wƖ�id�4B���0�@T`�ȍ4�yL�P�ö{d�0D����$P�_���JT.�0����m<��������OsFG��|��I����H����x\�A�!53P_+�TnI�b�ˎVT���+�}�	�����jz��*mY:�s(E��a�nȋs�^�T3K��p��&��Y�D:���?����06�h7�*��K$Em�N�B�2�gγ��с���^δ��6�Sn`�����F�� �g��9}E�[q{z���r�7�Pّ��b@�@M��r��ϒ���k$�;>��fCi��6P�-�ػ�F|di��7>���Hտ�x��D�\��h��}+�2��w��t�{�5ҿp���W�T��8':�σm �L՚U"��sj��ýu�n�Q�v�/X׍D5�r�.���tu\�3�U��3�~~#3�=L�c�*,258ai�̰���s>|�N�ꐡ23;5q���F�1�k���<�fg�+n��=G�f\�$��^V#y�p�!��E��"a�K�?���
���@��d��2c�.���s5�e�	8�3��;M�BpGMJ�2|��ժ��sX�7F�X�������Uʹ�P^�|!Y���)4i��I`������kV1}e���EA.o�����ë{�H��ƃc��N=�2�c��{
/�~�����5'�f%p+����ͳP_�V(�Y��`C�vżl�%�]����]���>T�e�����!��7���`ɫ�}՛��D�v��ʐf���ȸ��-��_{mf:P�{�Y42905Ҭ?�B�s݉L��vQSb/:X��0���}��Yq����mL��� �81h�����GplEL����Aj}T����oM�ƿ `(�3�h�f6�"DZ���K��=��4�ȸ��T��#�v�	��v)��"3���
�Q�˩p¾�ʖfK��.ǍS"��]�5W
����:���_��	�5"���Hb��Ȋ<�d�K�˚˼&x���jS�D�^Z��r����D�$������.	���ҩ<y���5�Q��,�a#W�w����t��2���5�� I���.G�ZzP�l��
Q�����:	䴆��*�w�,f5i;�&
n�[s�HʁIK��-$-�vG�/�sm�a56VO�E\+�K��]�k���-&j����ӿƅ{�Lg�V�!�q�t�� 3&ÕB�>f��dC#>�4?T�ȣ���'Ȫ\u��9���6/�A?�� ��s� 	�
W��-�l�ʇ��p ��2ح"�/_3D{�_7 x�`�s��#�#D��ZJ$�kF\�b\�ѐVF��b����#=g��,��4g��v��4�^m�pl�U��$���gW��*�R[�K@�
�bp�6�� ��n��{ph!� Ar=6}�}yƣ���}�(>�1�=��̵��o�'��L�4�D)��g"P�(=�ij L�*Jf� �ūǵ%�g���i�m	����}V� HP�8p�����-*F0Z�$0��TS��+��(��g���'�e=L�WUX�>�W�ה�:K1#6��O�]I���A�ƇX
��VBu�s��ŉ�콴��5�u�!��Օ���@�Ŋ�-�Kگ�z���uۮ�z��g��\T:~��}H{�y�PHL�H��}����������;fC�D�_��"%�7�i�߃_B=o���̹�-�� w]T�t����K	�O�ʩ�7\ۈpŶ�~H�������o�vH���)
D{Ab8
o��
BJ�J�v�}>�}B:�Aߤ'$�X.�N"���0"ㅣ_���_=!r�����s�忯ߘ�N��n~x�3���&P�Zt�d�TJ/16#�k�5�􁰞M�%�q8��k��˘��c�3�а_s
<�LX���}>{ӵY�@ �k1_�l�ȃ3���u-��A�P='�T��cgxe2m˂{T�4
v�s���LJݰ�#S��D%��q�q�'p7��2U��(�R�a"����0^f��og��i��f7����9\٨!v�g�Vi0��"I@ډ֬�4��v�N���ON�7�˒�	��ӅQ"�=<�JPa�Nq�Ki��b,�ff�3�\�O(���2��eڞ2Fk�#8�D��4��ߍ�-�T)��^i.}VV]�%WȲ��`��i�]�O�:��t.�;KM���lgHa��]���[U6�@ڗ��\�*<�	sM� ~��v�R��5�Ϸ��#d�/>�ާ/^F\5+h�p��L5`��W���޹��n���,��b��y�#vДSZ�PYo��eL����V��1 j�س�����A'U���.r"dR�-��X��x�_����:n.�Z��w,��7εjx��
�<��[�;���Km{���yz�����,o[�e���1���f ?BJ��l��Uxe|,˪�,���w��fl�w-�]���'�����{D�M)'�����Н�A4���J���n� �N��E�D�ۉ�eh�'�a >b�p���F������e��I�>�l\ H}���w'	eq�;�@����t6l��v>�+�Ux�R�		�JlK�,�J�ۂB��f� �x��
&y'b4f��ܜ�;W���]���m1|-��dK���0�cn7�Sa����u��+ 9�o	��`�%����Y�Y�"�4���>������UрNS.��1���&%?��� ��y�U����^�1=�om� Z��	Җ�8/ųĞ���1bp$b*�&�Dʝ!ҝ �������'��y$FWEĥ<�^��1�P4̾tu��C��m8P-��L�a!5y��f��ɏ�if������L!�8.��n�j}`�����E�)��v��x1q�������Ǽ�J�=D�kB�M���8�� E���p�T
�����e�ߚt�!Bq����ƿ�(s�:܋��.���Җ�1�;�|�[%���n�0��;?o_l3�Z�G��]�����y`
�d��{�Sf<ꔺ��=+Ǚ=It��⎖���h^l.���S��0V�g���|�,ja�է����3��O��z}Q�.tN�ms�1U}����@џ�E]����r����m���Z|�W��T/�>%���BQI�X��ܬ
�@�:$���W�o�XE�,��u<�9���r��ל�����P�9M��.��P���l%�I���� Z��odVJ����
>��4�JF��[�҉t^��
צg�g4�2���O���WDR��z�5AjS�n,�C�
y��ڦm�޲}^�jJ�Q������wh���ic���i�9F;6K��;u�+�Թ2����\�>���U�����'Z9G��f>���!�8��~x�AA�u�ybHqR��FK���G���2���#�M�b�:"������ڙ��b�T.�T��6���y]鐶f�>��������{����$�r�2�u�~TZ��6h�)7b7�R�Z,�λ��}���Y,x�Ңr�闯�*T�N6�>�J��뫖��_��zu�hK�3����];Ǡ
Taf ��zr��u�E�}	�'3E��"����;��ago������O{�Bt��J��n�~aڝJ���Y����L�eB��S$~��� >��>��O���:Y*h���\��եVy$q�a	ᬞ��J���3���=��V���ݡU|�tE�� �"e��Y�{�: ���Ш��A9>�7=s�ْ������X���s����{�ʷq�d+,�{� �b\dV�Fl����ok.�>l�9�I�4iWX��j�F
kn޼��
W]����O�Fs��Ö�u��7V-�jN^F�����A�B���?B��/'>�1|������A=���[�=�����[Bt9�8�{��g�:5<8Y7kU�]yοCn�� ?���QOt���#&�$��x^��kg�x�J<��s%M½(������Cc|4�����k�h���f�2`�L�QW�-��uT�.dBF������F������ڎ��8<베ά�m�gT�J����I��+ �#I���^D��v�~%z9S��Q�Xt̾�-+����=�^k���ߤ
/���éW�;l,T�q,��%E�s}C4Ԡ�Ng�8��{�]�:|��/�����'y�^@<(�F�eu-X"e��Z���M���-�P���PM��VY��Ϝ��/k� ��'H� �b;6�G�7��P;5��@ �'$0,�D�����R�N�<*+�AE&��ʹ�s�,��ye´ŝϓp����o�K0��������!�C��bz� u�`���R���9D�U���]�Øb�YږI�S)����U��Ɲ��^U���1τ6d�R�M��`���_О�}.!��{(���� ���!��[�{c]�)?\żn%�-Ϧ��9�K��?UE�Q�ۛ�|���(�ܴ��َ	Ƭ5�JL�>,�����%�jc��Sͳ�]K�U� ����
��r[@��$ט��i� *�D?���`�وq��aGy�"���^��)uW�"� �
� 7_q/�M���ɬJ���Cx3��Gk���p��|�,��N�=�vS�':=�њ̾���t�y��q`��2x񄌚� �Zk�'�{�≓�>��a�n[�wl5o}�ʥe͇ɫ�kj��?��B���ٚ�՟�Lcl�}	"�j&�'#Yp{KSu�a�k��*>�L��9�V�X�1�l"��L���=��� ^��/�K|�O�R�J�3�C	��#f���ZPW�첲�t��A���@��i��Zl"uH�mK��-��k��ϖ��ЌK�"
��M�@�[9-�B�e����ӠHLv���0��qzQ��4G8�+�..�O�p���kk/�w��NsvY �R镳A�?�<S����ʸnR�wť�#9�4����Nř��eG��lё�B�ǯ��.N��C�&���>��y��T�ncgcʝ��rq��sk��3~m�A�z�:M]]�D���T�'z�4��m<�ܡW)�T�������s����<V����Y��ɋ�O?�堥zA�25���7��Tد���-EQD�|���M�o��$�}��O��� 9L�`�y�b���%�� �qm;��=���x6����c�n�����u�]I�{���m̩�-gָw�dv/1~����wy��s,��J�A�ap���'��gR��DKF��`���]O�G*5N�=�^���8�3&}��_X��y�2��;�!���އ�~d�f��{d�H󆇉��=^�ǿd���	7t��z+���r��24����M�nIO�:	���A ��]Җ"���8'��Y. �r��]{��Ki.�`�K�Z8���~�b�g�q��YH�л�Ш��\Q"Ib��A�<���y�h���9>w�tX-"���Y.yPJm�O��3��Qͯz`'�v�:�x���h����g@&��+>ҩ^�HۋuJ"���m�_��#��4ȁ�)\,�'��#��⸥��>T��i�٥��枠�81�ԡ!��||2�C�?�_M/�:����Ri���?����g�wm�_G���Ţ�͈�� X_�x���֛nl�Ά�.9z���O�M�±{:��:�y��o�,� 5��AE�F?�	$�:�ͮ���1+Wg�Ho�`��izw���_.-�w��,vq#��G��鹠�E�Åj��qH=�0bU��\E���p���h����}c�YM��O��	P��ڛ�N��#��+��hud�M2�k�{��O�����Л ���
!"A3�#�	u�$W��5��-:x:�l7L2�R��!�j��c�܍��.U�A�µk��R=*S�P�`��FL�r���߷�t(����e��4m��h9ķ�O�FGhZ�V��H����
ߎ�V猑%e��qAKޯ|���p�HxD��ǈ�j��\#Tջ���.;��`�Y�.��$8 �0�Ƞ}~ĈN3�I�Lڜ"
�����w�֬���
)��)+���5P�jd?AE8zCD�d,�&����6�^�"+�^Z��S� 1���[�o�y�gz���1B=���Ck���y%���+^��w���@����X!�٫ht���W%�C-�w{��璹�p�+�yb.N#���S��Rt�h!4w@xww��},��̷2�[�jT�1����=>� b��63�P���P�q.���#02��O���;�����������¶���禾�Aa�Į��r�j@��4EEu�y�oi��`
{P"d�Oro�ο��w{2������S����T�w��Ż�[�A���������Srr�%��=k)� Ρ������k��D�Ï�vL0ŋ��{�%1���*���-o��O18���>�d��D�s;Gdv� �s���o��X��&5ݏ���BU�ԓ+�ӳ/�sñ�	+���:`��a��i�j=w�mo�>RW�J�q6Mk��m������9�� �Ic�UR�:&�{,f�<��7�f%(�t�
�{ff\����LSg���nGW)��,�KW�@��*V'Q�ǫ����Ƣ��(\߾Gb�����X����\���~A {�f���D��×�*B��K��n����S3�Yav�k�K����Q�(b�ĵ��a#���,^((�z��#U��%�I?���J�#lR�f�rX�o�
d�CUp_;����;݆���5��Q�|�yQ3�-����Y�`m�,jN��T�I�>C�.���C�t���x3�4O]E"��K/a�yH'oܯ��7�Ѧ_��rgSoߊ�8����_��D�  ~c�{l�0?�Md���Ѻc �ɒ��+�;P���Zv�����Ys"���X�ha�e>~R[�a(g��'q�i���c�#I)�~��B�T���b ��5�-y���Ȭ�ȓb���Z�SK�d�y�7٤TA�[Ι��}���Y:Ô1sbT���𧘿җbW�kw�ƙ�"�,���"�����ʾWrxƛ`�+R���>r�ʒ�D���-��tZ�ݙ�Dշ�m@��'J�t˽Ae����|�v�� N��H�t?��G�)����E ��b{c�eyC�ЧRY����s2�?��Gv�^'#�E���2J���a�V����"@I��,�5�����q��@k����!C�q�Y�E��x����?w{R@�{� $\��{R��I�����}�$�g{���7��f`	�ۊk
P�I����.֭v.\l:�a|��ߘ?��u�d�z����kx9�	7D/E�����W���Ԗ�oXO��AD��V�D.����Vx�Kï��k_�Oν�F+�$��>�,s�:���}>[�D��)�L׈0W�^V��G�O8����ݧ��3���?���Y��j�o���ɾ�u�K*��U�7�	܈o'�6I�\v�����@?5E�����I�Hghho��"[��lZ)� \y�>�$�Շ�#�{���)C[e��2��΢*�f�)L7h�G_6h1�I斫c�.�&����p}�|���=�7=O����
3j9p��q�A�U�&��g�2Ҧ)�**�C.D,�;�?��Ys�� ?��2þ�����/Lh1�O��>K���; R_����
f<�-�ߢ�;���~�>�_<��d!@�_8!gոpz�\e8�F3�ܨ�㽿���qbua�оq`�T�GE=j�8䶤��/�L%�k�%7S��B'�,����E�:Eo��~��:l9/ή�J���B��z�ݙ�!q\j����2	��S�Q���v�����w*Ǧ6O��=A*���1yi5���uGs�~m�EG��$1�*0�!XGLk�6,��~7*\W�-��8Z���J�{%!��~��(j���ќ�� S�qo�p����/�ݽ��"��}�R���L�y=V�h�5т��ׯo�UP�4~�z�H�+���\X��&��N�Jӑ���f�L�d�-���sp���5g��h�p��d��-d��� ��^i��F֐�0���L�),��]��r���"-+�!�<	>P��ų���ŷ{ަRG@"\	~./:�jx�CuQf�]н_�\����#bD�.���jE�Ji���by� ��D�kZ[����4�R�l�u����1nw�O��[�,t�cH"�(��G=���;�������ެ�¶UH݄��Gq����,��I��PA�/�^�0�%#%��g���"�j!;~���)��߉���8N�*���|y��u�C;�!�y��b.�|	o�ھ��p����3�B"��e	,��	�k^�!����˅+�Ƒ�\0�j����U�� �'6Bg�}�i�6C�e#P��E�2'��{��A�T�Fq~����=���k�?�u_!�@��it�n"��}��c�H�]ٜ��<�Oע?��2yy�Nà�F�J)[w�K�I�ނ	+���g+;� �$�j-�k7.'c����ڦWQ�զt�������!�c��9� -�%]����B � 09i��8���$:E=z��L8��#���h�𷸘+/�gм�C�~�éupR�j�.�u�Um��d� �o��&���#�k�=���qp��/t�t��Z�"	d� ��W*�U����څ��>��#���D��w��|�8mW<�=��/��':�����%1��"�e�RTIgPr�D���c���.�苻���ю��^���V`J!g`��˂MS��<��G���x�i���jp'i�����~�.���}<�`CsSy��ZVC��aK�:���1��fu�(����D:`��"MsƆ�(cr�6�\��"Ў`O.�(t$��@��t�w�hk�K�mfp�8�S:��5����޹#6�&�mw�т�h�����ws�9���ଥ�f5�g���Vq'�/�2�6� ��^���H���YD
�nؔO��ڵ!E d����"��bZ7v/�U������+��� v��TH�d�47i}>�N#��8���m3n����θ*#�U��j���p�t�����d 2(�N�݂.��* ֏wȆ�[�J"n�mt��	E�f�w�Bk�/wre�,�T�ҍg��OxY�������<|^#�^�̸ҋ����Ex/���������D���n��E�np�HuF��ѝօ~[��k�����1Y,bR��[d�:�MsX�\��_Q�ܤR���]smH`~�t9�Q'u23fkif���fhe}�>�eEZ����i��5�K�>���4`H��������A����k�P�x7���ڪ=�7�+zť�b�5�`�5�٩,W�n������Pm�hɒF�<�Ȩ�sa�"p�x��)i��?���˳T[ ���x`k�]d�w*z�#�7�����M>���p�SJ�T�'d��f�ZE^���ɳ�;�0El':.�$�!�2�Ms���l  �\{1&Q��\I{��l���$��J b\#ـVj�����dy��)��J��:	Af���%����-�v�E˦8��ڧ._���dk)�:�mkT��4~t��˦k��3Qy=��ӔT0
�/���L�^c���'�Ft|383Ep�#Y�q[�1��
�u���[��u�$	���=�N7ы���%3�;�(fm��'טVA��Y��A�}���K��a4}�Q'�Qq2��*�����9�,XX>&�]@ ����
�Csr�@>��_�+L�����DL)�9�ߟ�M����x�o���H�R���,Uf!gY�l���ž\�a�� Vb��Cź�[���/��bH��$����@D`�/��2ձ�Fs�;@��
uY>����	�J:�%X��>e/��<,�&�	��j06�&D^:M��ĩ%Jc��(�5Kg��K�r�H�Ç��N}8JK��`��b��Ĩ�ŷ'=�M��<w��A�H�BW>�@���
%���7Q/�$�:���\Ӿܽ��|�U����$�U�?�_������b9v�[�[#S�9���7&�g֓��g+�8(�*����5�r�B��@��-w;��("=4�
�)'��$1d� F��&6+n^}���<Ŀ����W�����Uh�w/���I��Zg_�Z[��Bo�}��CR�>1�'C�&{�5"ыU.�����Υ� ��x���b��	�m���u���Yu�ߗ��uv $6�{��H+L��n�|�d��:
Y��`]��:��~��)����ea��b6N��m*Z�6@����Iٖ������O�G�lg��)�9��*����8S��P8<��.����L�5N��qP@hp�&^�O�;��H�. +w��>�Gː�Wo5s�ja�W�EK������2�d�����qԭ����㹔��R�ڢ�tK�c�hEW� z�A~�K�.�����X�%�ֶRG�g���=%�����d4i�q�<�Y0����'��9���pGp;�tb4Ml<i��m�v��@���
o�bT9�T�>�41�M��ʣ	���0��2&����.�FI=�DfrFot��\������,O�䏅����#�U�*��~5��Н�'\��9\����O�p?+�I����wn_�%]�%	��ŀr����ʞ��/$��emt�)�����j�[P�5�-�i�b�kQ����ޭ�EN����s;X�=������+�����JkPք�6�cf�Q��C�u���fR���Ε�җ��lr��!�(�8b�N-&[蓜ݎ�T�T������_xds�i��u��ɞY�@4�ʁicO���0��W/�m��Wn�j���p�/�ӕ��I=�#k�����;��R�c ��͊A���4l+��3�e5`pe��79G��;N������&���o�*��8�0�CB�5�p���~�oZ�z2Tcf�r�����R���w�u�#�L��E�p���[Ih3"�}��dk�!c2Wo~tV�q�!>�I9�VI+��������Nz�x�VG��#� P�ޏۙR����g��`b����[����F}���>o�%o�Ώ����7%�$'���q[>��CàD+�MQmOU���H���&��̰[�Лx�)j�V0"�j9\�-��(�X-��q�ZD�H(�e�8}�
lo7�5���!m�^Ȝh,�q[�N��x�`�+Z�O���\�W�׮�jty���e��U��Ca�S��R��@%�NN!*+��d�-<qϙ#�$/DX���n12�geL#4QOt��M�C�.�ObB�\p����6���=`D����s6�� k���q:��2�m��>Q�?��|� *��������;��J�]),�����K�H�%�u�!N�𲛈j}8\/�l�Z�$��J\�<c�='ebo� z��{�%��Pu?\�{"�(h��:�E�"vPP�^v��63��^N��84-T���a�`qwd&�P�eL�p���}�\����#���Y�zC5y \�^f,lYu}���F'6���Γoh���K�D�d����'�=>5u]x(5�r��:��MdߕRLh
���گԐEt]h���]�^��h�`-Y�3���@�^�>E����%�|��<l5����
F�ΙԑR�Q� #~���oj�#[����:�,��R���V�B:}�4L� x���$�%��N[J�t��ߋ�u~ݻ>��=�/��:�����O��S���.�)��'p}v����PH;*�k���.5���H�oB�� d@R��=��(��*��j��Ji�]E�Q�T���(A�+�d�>���9�N.�,x�95�g����T-�nr;��ʗ�XR`Q��{v�}ۻ%�_�,}l?��#�R؞
T�߮7���`3&����Ͻ	Υ%��>�'�x��Ċ����fF�O��-{���AQ[����Ô�L���F�=[^?�0y�m�����B(~ ��#�A��J4�6xv9B��}���^����g"��K���GB�V��K�2�,���D����8C�'j<����<���v����%ǧo�MS�Gv�+��0��h�릪�d4�'g�#b�w4x^��eO���yЪ#�1��C�m�[������]��G�,�P�U���~�X� ݢ�;������A�3���z��ė"������ �)�m]\]��yDu�~ ��-P�/LaY�T�:đ.�e4��☆�a�9�����g�j�]M�:?��J�aЮ��٪�?۹޳ZZ���٩�w��U-���`1�tJx'�#q~-t+io�lȺ�f=2,U8.Z�N\�1x��h�b����7>+3p�Vc�3�9��j�-��o�3�J�q��%Vғ�~�q����d.�	A���L�{�iwɰC{�3^-u�p�� �_�[�CuMC��Pa���8�$oԜ���'�����L���-"�XF;u��?%e�O)hD���� S@�����5��i�X�����ll��Φ���b���%%�O�a�ˢ�3mi�<�d�M-ٻR[���"rw1�4D9rOF���vs�8�;�xc3$��+("�e�ۿ���sB��LiN�ѳÝ��|˕&N1�]'�=q�� /i�WSD.+��#���H��,n�`J�v.-w�٘�^��J��q1٘�rx:2�0��ɠ*��o�6�f���JF&��P��8����<s@�����":}��6��p�5��q֤��g�h�*$qb^�V:&J�;�"�M��������3�V��n;�ʱ-�T��3y�C�KY���BnTcFq��/�UE�����\H>��_��Y�cF?��)@Շ&|������A:��	<�D#�t*�d�3�����J�%'���A�tÈR&I&��6�}n}ĸ��_�߲�O��d �o�Cr�9����ԘP���5�"�!s3�Õȵ��Cj��OnW,T�W�9��;g�͋�+�96�Ѿ]�#�{*K!������y<���=�!ӊ�Ҧ��8뢽}uT2�b�+����ب7��$S���Q�q�b��������Ç+�1*h�)g��b�$�x�%��F\"��^��P�+�J��^��i��1n3�V�=Qn*ȋP��u�n�`j�﷑�[}G|�X�/1�n��K��X����Q��,��t��cӞm��OB���0�BwO�[߱�뙭4U�4�.��+�iD��
��0�xj�]��#@� @�(�� K � �}�=����
O��#^w�Fժ��f�7�ժ���Y�PY\!L_|�4�x�Fh:���C�g\n�*[��N�Z��\�qS���L�U!�s%��A㮝�s��Y�fM�W�ڵ��r����iZ����Q\�����ɺ=�0�SQ��%��W��0�/�����a
"�.�M8zh�[gP�,o���5rd:H�g�7�Ŵ-�R3A±ӯ�ik94��,ױQ�(�)z�,����l�+�3J����,���ɝ�����4*<H.�6��l�{]]r�E �~����*M�x�B�Z�+�}E �R&�����hS$8�š��Q���2�	P0 xj���&W���!=�q=l�i7A��*x8񑑔�.���ӠG	�)ꔍ�X������:�۸����6�5j0H��� ��.�|	����6�1��!�����	�צ>�7��7�D�[k�]te���"�����=���A
�"@f��T\GPRo��_=8��)F(ꕌ׼{�7O~�qQ�@dQ� ��"M{iFyݔ��	\����@L�2�4VR���u�`wY��7:�9�D��@�i8,�&���h	�?�91%�j�#3 !�W+���%�8���!?=E,r�b�>rm�"Q��f^k.��S���y�Fk� M�%@~�k���%�bǋ�h�\?�}q�
#�]KcQ�3~�6<�4c�ͪ���
�DR��U�%��܄��=#��3�M��6�r�̄[T{�������D���Op�;���U��X��qb���������$��8>D�_�2�qeH5PO��������~���9M�0ſ�^����IB�U�X���ʹ�э|T�-���5�B�^Ʀ�D_������)��h4��mf<�2�Ihv�Ʒ=�&Ѡ!�.>-�֎�@軒q���3�%��q�T���Ig�DP��� zH$�#�>&0Lگ����Y�#D	Ca���@��w U㈖�h�x��`"a�Y6I�����_�o.�`�,hK��w�AX����%gwZ����g;�^��ڥ!%��軪.��%>��䳏-���H�Б�S��OZ�oxw��m��v7����ٸWt�/��v5�@-��]�L�GP��4��&hC�8:r���kߢ��zi+� �Q��]�&q=6�x�tۑT��&�FfP�`$����!�N�D���`�w6�ﬥPA,svWt�j�Ƈ�o�d~�(��U٣ &�̈́�h� ��j����Ӂʢ�,! w>����U02?���>@I>�H7~��Ԍ+��^TՓD���:b!%��2�X���8��2�FY`�n�1E����n2 &T���c�jKϘJH �p���~0����'~��a-�PH���z�w����Q��4�*�LW7#��FG7O?`
 �<�-���yK�����~#w���|�p���%����v�ӏK'�͝�ȥZ�n_�WY�j��%�[���,&�y����rZP��Aj��?�Y�PG��a�>`ZK�_�L�1Q�u�`>�ƃT��:O��nq #1"b�b�e����$Rk�>���9s~�$�� y���r7�ؚu��r+s�Gx��3e�����:�����>��m��H�A�dq$����oJ���h�lT�1�����.�V˳-��L���ce���^EǊ-���2Zm�x�ɸg=�,ac� a܌4@���h���ZI���:^�,�'�Q1�B �����w�1D
y��b��I�����V����T�T>����������~x��\rL#��AB�	̍��wjJI�Pɸ��u�J,����v���n6%��%;����2E��33[�S�.�'@.�2%��l�gt�R�Bg)S�sK��E���J<��w�ʉ�v[s@$A��ne�6U�}0��m[ZeQ&,���8`n�J�������"/&,:X�ov/%�� ��<���ӏe��+��_Vt+;N��1)�҆�mms�?}�-�v�\��O��%��6���O䵚�0�=�ܫHs��e�)PA�� ��z_\���s�&���&��?Ns;�A!EL�k��\����з��9��&�A0�
��V�"i:��Vq���\�jB�}[�Z�p�h��{�iw�f�#.��H#�mWn:��ع��L�������_�6�[���i��S:o/
P97U������$�6#��jT,������X���)Ю����S6i����Ϭ?��Z�a�QWv�0���
&�<����Uj��~��l��(���7Ь9eh;iORDϹ!0fR�.�X�mOJ���Ә������jo��q_��� ��|S������ZjZ+Lb%�rڽ�f�����\C�5����U�վZi�ɵB�vۊEE6�����4ќ���1"鍞2Z��� ��0��8P�<&��,�_BEnYe�����ARݝ��^ǿ:N�}6AX����%B��������Y,\:%�y���Uj��5���Ϣ�kg~��K�p�~p0^n��c+����	Z3m�-�y�x��'�Ջ�h�e��C�
,Ϣ����W}�2��TDԛ�/̚,FCp@�&C�?!������x*���}Luk-ŉ�<t�1��_�����~Yl=h䝂X ���U�e1��6���4�x% ��d���)�{��%K��_��,*WO���	������*�F'S��k� �tId�dR�����"�P]y<s�b�C#:�Ǜ9j��������{�[G��wᒸ�AQ9�*I M���Î!�p��Mu�[�pp�fhuht����^�O��:�Bv�����������d��~`.��"��E:r�2��.��sM�\&�¿KF���5T�>�!��ljx���wx7�s�x�-��x潱ty�	�b���G��8MO�'J���7�i
�����7���&��)����Ћǒ�=KEÜ|�(�S$)������cs���B�����(n�	�	��3��ד�A��������J�b�19D�y�c�	q��Z���`�U��eS��s�2��׍2{�z5آr��n7p�lyr$6v��ֈ�Au܊�w_ՙ>��c��CX�֦�y�����ܓ]?���0�YK���B:TY�BE�İ�6^_Ւ7��mw���/���,(i�N�`�;0/ץ!�Y�CR�fj*rd�K����w:�UU �R�m@h���O#~o���3�
{7��-K�n�r�X�p�e�њ��P���{0�}�ɣ=M���K��B_�U��z�{y�(+�aD�Itc������������>T�\ �� �d6g�U��u�����2�
��|�ŤE���ZM����6�3]�H��C"Dx�|�9Є|T���Z^71S�1��x��Z��ML�d�)*ޫ�|0���X�D)R�ZI�� f������s�n�����:f�t�.S#0�4ex���ە����:Ӥ	�沟�̳�Ң\1�m��9��ih�����]���ɾ����HM~��.�w�3iO�|F��8L�8�+����d���!
�p1@����F�]��錐' \HMfR�Т�s�,P}���IJ�v���lCӢ$Rg}�҃�Ç睼�f�{t�3p�i�&w,s'�����F��J����I)��ٮlٍ�y�t�c��:e�RI�(f��h�Rø�0�fT.�-��0�*:�=e��U��3!�g�`u�[2~w�g��:�0h����v�yb"�|������ �@|���{�&��X �?S� �D��x:U�8��G�fDR�4���
E�I�����zU�W�� ��{	E��{�O9�h	H�(�@��!�^���Di�#�螤m��]�o#% �U>��K������M
������� ��1��đЪre�����h;�
����G�%���ZP��CgBg��D�e b;�m8i���L~ZT�1������8�\�Ds-�~��Hc$Vp���3i �z23���|=U�x9�[�ن��������-��Lq � �MDԪ�[�k�����86��t/4�rնYN7���xF7�u��7`�	B�nO��} H��R�+�/!oUb�ð6�{RW�}�B۾���s�Q[���(a�//lT�㠯<k�ݑ����'D'Lgc��y��W_ ?�:��/��?��0�e�I�eY����7�nXQUL�g����Z�mjG?$YKk�d��s*W���pj0��� Zd`�Lt&)q���̎��Ku{�{r�>�W^�b�,����l�M��#M;P�2b������K�[�c�p���,"Z�v�ey��77��'b��Y�����i�-��$'E���f�)pY�P$W��PJ8�3����Wj@W��E,A�7�vq׃Y��Y��,&������KW���ܑH���ǟ ��V��geuU�)��1̴�}�wd��Ny��ʢ�fCt B���'@8��4�N�ƻ9%=&�~��0��ճ���Vk�@P����3��Vb|OD�Q)���Yf��@���W�"o,͞��iy�ٵ���a1���>'�!����Y��_J��Ko�5:f>����Y/��}V�#C��$iЈ�
H�����.����&���K�Z�+�O ����p#oq�pw2����Щ6����N�l�o8�� ���a]�d|(D�7��
���ArK2�E����#"�@J/��*�1J����w�x	�!��Vŷ���IMЬý9=�݀z�5x&|9h8Cǅ���;���*I�y���	�6��%����Ȭ-Ϧ���u"���#s�DϸY�.WFЯ~ʚ>�\F����9��].������Y��¶-zoo��[���4�"�]:[�r���;wz��5�ҩWpy�J��ʣ��B"	zN3g�$���xv7Ұ|qU��m{��� �n�����$!��K(���x��W�ڎ�)����o�|Q���`�{�$�����"��}���0O#rSe���d�3(v39��̼���6�8��l.���n��)	�r�Ǧ�W�;1�=gB��?�@�З�ofR�*�:�����h�m�<��%�n��T���k~�B�S)h�Û�	�^�"6�"�CB&�m��9s����l��� ���LLg�� {H����e��t��F���°���M�Ɔ@5w�щ~��)ԗ��m���ᗳj��oӦ�ƌ$��Gn�C|��p��d>c��V����s�]���*;�X�Ur�lc�҆0��z�pDT�������p0r���
LЇcY�h��>�m
Р������X�����������4p_'�Y�o�xh;�j:[y����������Dw����m8����qYD?D^ܠo%��N���J���+�E�5�X񀋀�1�ʀޯ4A�݋eۿ�i�W�x &�+��R�p�H��!,�����X��:*g��vs��I�	t�GHV�B�	"|g����B�?G�x R����E6���$��r�|��q���?��9��Q4f�?C�MM(>��a@3���V�6W�ѳx�*�3w�KHS�1����"w�e+�6���t �H�N-�Pe%or}�a�khy�=�B���8�8L���q�E9ݘ�+ρ�m���v�h�tՕ��sۿ�.%�t��[�C�w�ɹ>��{0۫������]utx}�A�O�(%=�E1\�>�^sv�'TJ�����Gm������]�J�S�S���|���D����p��&��էLCl�*�;��I��$��#�m!1�l΄\C LW��Pn��+�_��ӵ����'�P��HꔧTܥD��B7���(\�����#h�m���Ps2��C4�f�v�U=��4�&V�4��aD�z��\6F�=�nm�6<+�@�/P6��iX�����>NZ��l[M_l=��"!�����۩����P>�d����JV��3�G�7��o|�D���ԩ�U9H&P&�5G�Z]ϴ]߅1���������[�e2�aY�.GE�����"�:\�)�G���XD��Wa?D�� ���QУ�#Ffg/�Eb0r�	��0Y �������,���yZ��!@���V$bN,��6%܋zQJ�J#��Gg+P����TY�VզB��#��!��%�q�v8(�7�BtI���BN�f�Q��[�Z=�]�Q��<��`$[�k��3�G�އ(��7�Nu�����Ԑ�e�W,W�^I �]��f���%��|a(i�H���S*x��A��3�lWU�A_��y��S炭yS��]���TP��jq�H����;�YqH��&��_�/Q4%�l�̥$�D+��-���D�n��͢��d�a'�U�A��g+i�\꤈c	�b���J�UUl�f\<eFr��SY��<�Q�~߸.�����7 ��~.H�a	p�kB�Ȕ����N���k�/TIM�6~Y� )Ύ"��-�}�?�{|�$TL��T�������=��z�:��X7�df�d�i��i�;ή%Ȗ�7+o F	�-��۲���~�n�j�Y�aY������5&rw�F�7� '��L�?6�E[?aV�EG��邎�ƥ<cNnq{(����{��E4�cˏ���4��i�#�h�=y5��,ka<l�p4�yU*G��*�	�8z��T���#�L�i^��r�����6x`�]�aR�n���e�*D�DP�V
��N�6�c�h
�u\ [�
Y�t7�T/*� y�@���7w���W��<d[� ��M��̌���Txl���3��"��r3��X��u�g#�S��0t+�W/�/�4���5gʹ�^��Π/��B?X8�*CS�\Q.�k�<>��hO#��!R�nʯ�eQj��@�`
ݹ���iM)���5�S��g����t�A^$�drƃuI$�[�!�^3Yd�Z3��S��Pj��6@�/_��wF����cr2��>Ӻ")��j���Lc���1���ٽ 0��q�Ԩ�I$�}�!��N(����^3'�Ä�.��ʾIO1+\TlY�;&�@G��oD������H`-˸2�e�$Kuo��Ŏ������,f��SR{2�4�̃M���[�=T�(p�dO�')�^1�Mֻ���(�Ǩ(yw
l���Gd;/p��q]]�MLJz�pȚ��R�02�1����`�Z���F�0݄���������p?}'�v�?�#?k�dWI�/��a��x��@��m��u'�)��q"^L�����/[�f�^u�E���-��>��	44L8v�[a�uߦ�6al�J�7U��JK$���� �\���V��*?�'Ӯ]s�&~��=�%1;�s3:�j�WE��q�J�����`��}��L�Ӧ2�=�~�2�����i9����Z�_��2�YhW��-n�����Y� ��7D��-a�0�C#6�Yۦ��U�.��_��q����Wt�S�3�}����-4�3!��R�����=)c�h�xRB�U�F���x|��8�J�j>���
m��$$�]��Z+#eћ,�t^F��&֑�0��M丹a��1+*�^_ѝ:��K^�a���ǧ/�Z�fW���Y0!&$�x�k�������C�}8�b�pM	�{ђ��&8�۷7���9��zM9��v�Q�N�������	������K��Y3>G..k-���kfR^J�/�y��Of�#*��*�mw�7h���\�i2\(�D�E�aZ��^��=�M������d3�l�05)�	V��Q�~��Z�6�ut)�[��>��n'���M��xy�66� ��tF����5=v(Tǚ��f�g���� ��2ٲ��T�l�[�g$���Q��a줍!Er
f	�:eC^���,y1}k<��������7H:y;��uuQ�:�<�X(��9#��҉
\o�\����a5ʦ�5���n9%hX�S��/������)��I 8�4�ֻ_���#��u���&vG�Ʊ��S�(�Q��D	#.�JD��b�}>}<\�� �8�g��s +*����kB��n�d�@;��/��[�M䢞���PI6l�U�n@��VM �L��ݖߐ��7����q-�Xm�3t\�j�rm�h���ڡy{o�e��&����:8����p���3zI�K`��� !��3��,�\�#z�@�gW`\�~&u�71n�b��8�Ww+g"�� �t�`ͫb!�m��%�x�~2UBU���I��xp]�
~�(�����-)� ^x;�"�����w�&(��V�s:A}أ��u��Y~HqG�T[(K�}Xɤ��z-�>ϡ��/b��|;&��Z�������R��Pn(zg�ewlg3e��%��iNқa=xhN�FPۿ�]���6|cɭ�\���1�Wr�x�=ȶܖ�v&�(�ͨb�nw_�X��q����[��R��?,l��L:��}O7ŎbE�4º������B<�
�S�D}3��;�(�K������Jw�2&���g�,���13
E��2b�i�����*����V����
"�mط|�-�/h_�p�> .���M
Yb�B��MI��mx���F4R���@4e%�����T��d��DQ��Ӥ'�	*��|�jB�44�~��8�<�8��1AZf���k�f���h�H�`յ����5N����棰p�2q2�6$Q���?F�s����rhN��W�&�.ũr-����,W���d6.������Z�e�k���|������F'ǽ����u�S�} ���OR�Ha�}=���a���N�\���Z��`SGׂQ�V�M�f#�������[��ډG�̳'��6��-d;���Zw'�_K��������+5-T�F����T���R�V��JQA�a���)CC�Zd� ��O;�| �u-�	�����[���u���2͵wg+��	Ҥq�a���y���VR��F�+�F�(N����;aH�i�ӊa�V����������;�����p"MS�8��v�sF��tw���g�P���&�{&늜o�O�e���
����;�4"�j��\8x&�� �S�7������&Q�� ?ܮ��l~�I����(�5SN�e��*��u�+BQ��f�R� �n���=�^�tƍ�_�WV�<��S��p���2nJ^���zN&��N�%���'5\�}5FI����H?M0���@6g��b�w�G��G��YE�ߒ�z*�\�N�Q�t�Hz%ڨ����ä����r�'V��6��C�3}g��c^`��T���{s՘�5�q��c��LH�2�h]9+q6��duN:���_�� 
ͼ�k��F�^5�Y�*R�I�t.��aGW�Gp81�?(!��q~���+���c:<*!؜���"��[����N�;T�����2��������r'��Im/�zb��6�c�������Q0�)�=�
�N�Ќv��g�S�j�Ƭ�%�����Z�]
��a�����.���n7ι�B��>��~ΰj�8��O�7��msc��1yC��Y+��tG��h�'$�
�C
�ע���ug��BL7������]���`"��0�&_�f���W�I��}��o�Y.�dD�0F��#�c�áE�� �glG֣km4?�-A	�����a� �K�̾3?�~)	
������d���7U7���+��� �6�F^�&�a��2�&���cI��@O���)�����{��4�-@i�<�*�ړhW�x�*�z{�3��䛆�h^���o6���Lc�����3���Ɲ�k,?,8i�����iܽv`,h2XcņZC���e�0DŬ#+!����t���)���� �GJ�9�`ur	��Ot8��Q��P��O�9�d�)�w`jhs_a.o-�L���O7$��hxuOӠ�V�k����uU���] �g��<h;pѐY�b�����6F��d��P��8��Q��nz�g���ÛWOl�$(-��Z���~|�� TJ����$�L�ؿu���ےRC�\��:Z{������*5��
�m�B0��Ъ8�{K�#b^���ۢ�	�u�|�8j�������є�|�#��)E:hPr�o$[K��v���"��=S~���4�׀[90��2�k���,�.�i;�
Tѣ��G������S�	����n����mybb����q�\x��藺�dwu�?�с+�JO_q'���<���J��[�A���A�X�)/[|<����y�i�q�ܝ�������*���ͳ{5�w��9z��	�g�@{l��dz�Hp��,�D/�n��^��bu�YZ�?�z�P�*��FU�������tuY��_��yJK~���l=$(ˬ̈́�u���D18B~�XWy�1��<X�9�@�����u��)�`A'�dl�O�~c���@�>z�b�
�_�O(	�FĽ�j�K�[�G�vG�q*���'WR��B#J��?�7^r�w�����iOi�tn_dM��9L��{&#��{P����V��Us�����[�K�4��V�1�,� 0�E�D.�H:
����ZG,������$%�Da���G��T5��v�����(	�7������J��:��r\Fq��93%v�*��8���`�7]��ޝ�U�A���"
���p�cd�-��^�˹V,�hd<�Оq5u˹�f��[���i��z�S���y��AC�����������G;#7R����%5�e��˛�@�lR>��s��g	��C�0㎍�&&^����Q��,<0��m� �����y�V��^/0���t�L����2RU���<�9�	� k-�6G��Q4=��������P����a��R����Y��>��鏬/����E}~T=|�sVy�rA}t��r��:EK��2ߦ¹���R�rVަ�Q@Z;�8h��?׈;䷌��쟊�#������Rti���j:�[	��lw��5������֎5�h��/M��#�9��2.��sޯ���v��!��P�Dك� 2�e#�Kaa>�r�.('��Jw�.o!���yD �"c��x-��t,YyW�՗b�)}慡���:�y{�ʷ�c�I��]�<�Zw5���Fu��P���4��#��~N�d��|��s�F�l�χ\Z���s��X���������7V=�Z�K�t�Ӡߌ�|k�iO*{d6�������Ɔḵ��Z��vI�/x����{����ރЋ�)rP�gP�� �jϩ�f�'foߊҹ����Iv�"�a�=���*����8�R�t�����
.�a�3QDs��[����Q� ��܎G0�A�M=x���p~v�D�Mv�V�B8��X)#�4>	���f8`����{��e�=���n\����g�=�k9QF`L�Vu-�M�I���\�Qg���~1J� �xAד=쓭D�k�O͔=*w���1J�#E)��Z��;ğr�4��ϔ�NR��'8�)驶��τ3�;�=�?:��}Ŀ�9��k��8!��:�xD� -��|��U�9k��!���0�E8��j�7��`W;7z��Y�1L�Bx����&����Q�C_�x��榖��86̂�][޿���:�����zb���m�3�� 9��>�X�p�7c���v�~K���+��x7�n�v
'�ٽ��7ġ"Ӂ�ݠ�g�l�del�Ob��)�Y?zL���l�I${�����D2�ͱg*ω�*���M�rA���{
���AK���]TY�b�s���QI�@.���!�5��{$$kݏ�=?n�g@�\�=���m����WB�^~q�GN���R��K�Z+���	��	k-w@�Z�X,4B�P�l���U�'�-&�x&/��-�� = ��,Vl�1��6���)��d�h����T�ۊfhc���:���H�׬���NQ=�u�a^f�k���p9�Jq4]^J�٥��j\�����*ok&�yym�oB��vK&7��3�v�N�݆;�>4��wǓy�0p��@Hab&�AY����ם�3 �o^en~f5����a��C��#K��0���t��l���smܾd`/���M�5/��(o��m��h�B��	=����[e�� ���Wt�Q�--7Ei�N���oB��#�����
<�w�]J8FZ��w�?a
D��Ϛ����9��� �m@l1�1=7>��dy~���뵻����c���K���1�_t|���t����<��}�������D;`����u8����ޱ�����n���D�����î1h�jFP��:�$\M�DI��{4P�!�]��#`\�7H�� o�8H�/Ь�������F&l�;�ǾQT��߂�I&쯵�T7Ҵ���JK����Q���[������B�K��b��PC�W{ĥǡ'�aC�k�2��/��%#��-����v?{��T��c�q�U~�1�m�K�=�����q�	w��|�0�a/�k!F&.��v֡�����,X_vG�"��Z��p5l�R���_D9�1Z�Y�qHvT�&��3�>����9������C�M��n��g�*;I8��Ĥ��n$�G�ީ�q���Ͼ�t�r�<�RDv�u�Q�O��������	y�:�l�	�֯��6p`D%�x�Sӧ�Uձ��\�'R��XAeG�(�lEvUc�h��-!������Q�l�_�~��T X �Oާǲ�4I�8k_�ڒȎpc"Q<pnV�aM��7�Ǉ`y�N^�վ�]t��g.�Wd��Q��Ы���3��B.+�E%ѳ"�۲�L(d*w�ǈX��$���1?�э-R�ԛ1���q���������w7T�/H'3��o�S���NM�f\(�.����d���d�/��4�E����z�#ĸ��0  k�ɪ�Xb�=7�o�a���%�X�D���1u\�[dt"��ʍ���
3�kN�H��"P%�����y� ��(��	��)�P-��/��8���O�2��{����4���P/<��|���ԾG�����˷N<�Ψ�7YE�,�P�P;+�ࣤ~���v�E�$jM�w�Ro1	리F\����;yqM��XRj𯳼_7s�(mN�q�-c+����f��XR�j�p�8`A����_�3�W� �(���+0q�0�q��������yۜJ"����2Pb��WH"w��b�t�(�r�B�}���)�������K�"��z�=�����H(��"��%�ޥ�a���n�n_� �S�L�#,`�}�o�N�։P�f��Z�Ȟ���\TsTO4�v�{�6���@�x��*.4�<��@����	b'[m6<��y?���2���6Z�����<�."<�ӡ����[��Pϴ��('��8�mq�4�{�g��c��:ְ[��p?(
`@&w�S�.ڡ�-V�C �Pa��Z����<A��m��|�?��wiq�����Ѓ_Ʀ�T۰���"�M[u�k5����H���}�it$����K�y��S�<��K��]~˶q[?�e�����0lHH�fZ��b�����Ƙ�7�m�8��!�v�� ����)j�@��&����S2��؝Bw���lՖ��I���]:-Wq�O&^���3�nN'����
r~�6"7.YQU�CA4���"y,=�m�b�ҩE$Mz���0/�%\�y�*@�(�2�� �4��,�ˌ�+!{��M����h؃n��ȗ��h����9�>'F�#�����zF�hfSp*���"��M�q�L���i�9=s2�*Ύ�Ts��TcU���S�#O��"q���K�J͍�%V-ɘ�f�� f���~$c|��zGeH�y*�M��Mx<\��(��Ctь��Ն����G�8N�=�Հm=-d�ߓ���{�FH�L��//w���ۄ�7�ۺ��I�ҏ�^�.t��p�6���D�m����K�6�����:Ψg�Ff�%��7](�%E�ky���s,4}|�w���60g��b�;"���@�B��4�}nV����2�yVrB�d½9�}�(������#�착�pZ��H�NWC��D�s�)��k�E�N�0m�ϑ��%�U�=�D�}JODc�v*2,�g�֥��@��0�j��Oc�0�!6��T��喂�!���� �'#9�׶>��:�/��#����
���cՖ����Be���ז,xG_0��ȿ�r8P7oi3�b!To��蚙2,�a~k����y3��>����Խ������J Ej_"����o*MlD���/���5촗�	��-}!���l���=��	 �Fy�3��C�n�����q�X�G��n��(B$��Àx��#�����8b|�i�;
��Ɖ��f%��Q�)?��zo 7����0�b�\�W_0v��$nq�n��}~$���\�k� ��̟���΀ש~Fq�8��.�Ћ@����f�5A��L��2��s�j�V��{��-�P��{>m��Y�|�6�����C�C��(�E��<��|��g^������e��zO��ǁ��s}�aL��5nf�	���R#��Ѻ��{��deLw&�*�4�S�0/n��20�� ������tY�����b
6Q۟��B5���s�%�bn��M�=�����c�Sl��~�
�̀�̥!&YD9�:��ٜB-�~�6s#|m��KJd�b�bpU���B��֚3���{=��)Ϛ�A��r���`b�n�C��I�OIݵ���ջ5��"5�QǊ@:���r�����T&O7�֒*yk+T�A�{S�~²�d	f���ĺa���>=�"��MSå��-�v7<C�Z�#�]Z�ڀ~r[�)���O-#��h�{QG��#�C&��gT�o5t��м{~��x�05rM�#��E��I1����a�8�k��������ܻ����*�Aȡ���/dI�MϞ�*�ѭ��������]4V!�K�jk�G���2T�.�k��Sx�8���&]��4��P�^X�As�>4�7���%$B8�>��R��#�	h�"�x�ɍ�����0 =S�9�o���f���B��.~|�:QE�F��z���j��p�@��m���_CYy������h���8܇�Kq��t@��.[�W���D�q�sc�&��+�r�6�Z��`e�%��y9�n���)��'�X� ���{�wO"��e.���*�g���
|�p�q��'���*a��5)�р3�?���%I���=�)�T��G�Lc!�ï"�Q$3�73���g[6lB���`=��?��W��u������|������3����a�����;l5C~i���v�� �α�r��7�t���2-��l���4�@�u�]Z40�:+�p��o n`$*`�"���n[b�����*N��,��c�A:u�,j�e�z�~`l�<(;ϴ��=7�6�$�M®����Rh�����h���̀�#G��08�����k��`���$.�,��1�(Z#9��k�����7�֢��H:�85��Ǵ��O�g:M�{���|[m�%�v�� жX6��U~f�+|���)OD;��o���8��tq�j�߉��K����v�Jmr� )�SU�~�d���@�#A�k]i�o_oIF̉>��mL��T�6 ����ū�M��l;�s �.f3W��\�+��RC�~�I_A|g�lp&�qّ��O�"�(��ӠR;}�}(��MF� N0O&�>�;�[Tm�5+>��?��>�mϻM틭�/^!\;�L����R����>�̐h���%W����`�y�b��9zb0����i��x�2L֨�����ȃ�sۭ���f�/
�>��#u��MI��d0@�@����K�(��T���XK��&j"Hk�/}&���bfMC�F�#۽��渞�a�PF
I%�9?����` ߬+ޱ���_J�S�b=��L",gN=��@��:KB|�{��;��������}��0R�U�VԶFUew�� ZF>��6�f���(���ggL@��0̞;�+�`H.84�F�������Ѩ3����oQ�j� �qj)�9}� ���C	��c�M���9�L���aiBCFc^�p���;�0	��6V�Wp��=(�~`!
Ҵk+���zK}c�:-T�8V� ��w{�ʀ�
ڪi�&��čZ��ě��]X��H�?�]#�_�g��)[)�W
��0��໢�a�qWRX����ta<���$ټc�7�ݠq�V��P̯����Y�\1w�/�h�������dx�Cڒ���Ey�p>�#��C)ҙ��J�Ÿ���bQ�,�<��z�O%Z�C��*�k�+=`6�>y��a(��|�B�M��YT癅f>��]��
�S�D����|�_�p���	/�L��ն���ʀ�&7��$�m�E��@X��K$�3U��_1|h��w��}3�� ��uf�alU*�ۊ%�s�_�F��Q�4c�^Nޢ�>���83q�N�G�U���\���ٸ�Z_1SV�7���A�(��&�m ҧ[H��52Q�ܿ�9�|��5��QM!��swIC��9�X�l�`����vY��r,-�N�� ���0{=���&*��P�^�T������� B%:,M�p�0�h�ߡ{��j�93��8�AD�f�)ŖsT����i)�4tj'�:h�(t�N��65i��Kn�w��[|Yz�e,n�(����Qm���&��J���[�sᓍ��!�4,Y����?
rѥ=_C���͏�꿺���������ny�%�����3�O��X(k�0Z�pukve��!�8��G7uC�)f��,y���*�fRk�^��1%*�I���T��i-��z��
^�1�(�>���]�8"/�8��n2|F�j\���-e1g��q ���Y9Uص-,*��$�i�}Uh���4XkFRY0�$�y��K��X���c�ЖI���*�z��2�82�GU����ƒ���wbD���;��Q�S�
�Y�~���>�җ܇[s8ۄ���V�?<�q󏛷O�b���37�,��w����<j���`���3�i��F�9���|/wn�7i��py�S��G��5���پ�}ڌ;��Q,{R����@ˮ�8Z��%�I��79��iNn��V֋6J���a��k'�ce*��0hy$h򝘰���e��?�I��] $=�ȥ1�D�o�h��A�]L�W҄eh��ķ���	��dߔ����ag:��&�+�3A���/8���{�ҟ��ϧ�V�0�j0x�k���T�)1�r��� .��YVo	�tN"镦��|?�tE��C�z2��_{
���y�-�/o 5���'�Y��Ƀ|�B~�C��+@'�/G�!�|�1P��/;FB�{.�߇�R7�Ǹ������L���V�d��T;Q���gt,,�֔�ڡ�H�*� �2��Ϫ\iܿt������-Z|K,��L���@�J ��M����q�Ӷ8���S����� !X:}>�d��~@�Zc&�����6�cmκ	D�zP�u�E3�V��ި����A�q;Sm*a�x�� wش}s���	�90d\bM�]M�:�A�BW�O��#���W�v��B�:�f	���w�u�]t����}VY���1ׅi�C�|���q=#pJ���+�XhAw<��[ZB!�f/<}�z��^T�����\�/�,KS����y�"����Nxj	^r�\��	���y�S�QT{1yW
��[�G��q���\(o�O�{�}�#����po?uFy}���{Az�Ǚ��o�7���)Q�ٍ����
�f�;���}�y�<�zf��x�+��Ɖ�����}�D�Y=v�?��MK����8��Ay����R� �ُ�p��V;�5�B��&l}�>�t��C�U��Uz��f%����ۦ��4j³q9nY[��
{�G9��B�{�O�_v0�"��I���9�h6�j�rf���z��	��q�c��z�+��=�-WG��,V,m�n�{�$�؟;'�*쟛�qK'/�����,|Zq��/��3�
<D7Q�;)ԫ�u0a���_!���S�0�'{9�I�ieY�����[ TB<�r��PA}'�G�T�HQ�`�
x����YHϖ���Ѝw��u�/��va���|j�l_�n����@�\T�� ���L�������E9�&|������7�v0"v\��|=8>�!�����a@� ���:�"]�m$au$�N�(�����y��K�s��iBNL���3t���ؤ`��	%�Z�*hI4d��i�����KygR�I�/���U�� ��&e�GWqw���oF �[��C�G��#�%��w=���-fs-K�m��'���{� )�LX0��Lʁ���,c�yG��%O�q�J��.ŦR]��}s�����a�".��|�9M��Ҟ��~Ɋ�����f�w�Ho�LF9!��t�ͻ�w��G� �l:�¥ Lσ�мc�bH����<3vo�U2Wk6�7��)���9xsO�t�Z*��g�����w�i�e%��@���'��i0��d�!v���F�3�#�X�������p�N�Fz���{�88�ȗ�꧊�\͙�dKҀO1��Ë������O�s4s����#Y�I�!d�H��(98������$�:�%�*�{��x��e��E����959�H����U�7<��Hݥ��<� ���+9���^T5��S�D�b+�oa^mǘ���Rdܘ�۵�o�k���Q9V��_O��	ON�F���~�=�6��xKj�{Qa�4F?�H��wR�6�"!KD`�I�V�b�G�����M��٪]�� �z:O�=󈱣�"F�>�*g���bK����I$�n셢�G8W�>�i�d�h��g a�J''n�1�0n��8��b&��A@e�y����Vx��v�QsRېWL���e:h��/���A��V<�����ħ�+]�?<��jɯ��~�K���m?c�6�c�s�O����_��lk�44�j����,d�p@�e7��G�3?�P����f�j�Z.�-�^7딳��?�ώ>P_% ��E��g]gg�`�W��Y-K1G\�oL=��u��*��2��5�[G��_c�} �tRFȸw]/nF禤.�v{a�Qg���tҌ����t�ۖ$�R1	4�.�.j�4s��&�Ŀ�ZT�?���^���^�p�P��ݺdV/V��ڳY�h�v�J�ne�Z�t����!z- ���F�����YBk�q�-T�k򧫨:s�2P��Գ�3! i��sЭ@�W��2�X�o/Ұ<��e�߇�B�L�A5TaC�尼�@��ul��Pt�R�$� �x՘��z���z�2,���1Rw�o���5�m�Ϣ�%3يؾ��gO�l�<N#6P$���\�R~%�Q�8��m{w���1�2�cU�uP�6Gɥ���d�a)',t��|ϚSvG?suz�5�J�yRoJ���	��Hx]�����}��3<��C���G"����ae�8~�s$i<��Q��f������RE�^�>�r3��U�r�!'��Q�/t��~2����;,�������n���g[���s`P#��T�)�Ҝ�>f���$�ܿ��&�����GV����@�#���$}��c|�jg�&a>6>:�y�v��jR�������I����hpN���= H�7��{���"N�����>���RRe���WV�q0�b�iτ{�Za�ٛ�I"�@*ٰ*��,v�H��}��)J��"/)�n��9����� ��)�xm���.���ȓ������Bb�܏@������+�yP���=�}xt��m���q7�a�&�,�?���[y/m���G#`��]��qf�9�/>�|��uKH���>~��B��M7��y8�	+�1��<��ys�նz�1^��)�qŇ���d!� _$O�qT\aEŸ��S�ƛ�����Z_�ӎ���}����rց�QŌD�B�FCk>(����!$[�!@�"e ��%u�>��ų]�]� �7�j���:���c���J���L��=������k�~��c���4=^��|���7�y�>·�\�9;��9�߀��� ����`�pn>����lt���O8+7`��f1��0��Q���](�HO�Wi6^��@q/�k� �89�Z��x�Fa�:�oSV4���ߴ�d�L��/�������?E����8o��{9�Q��[���"���P��C�^!Y��� MBD!�N_���
]"a� -���.�kch�t`�J�%��dl�F�u%rK�iF(��J�I����&��5�
�l[��%�|�Zx˝&�/� ���mC�#T=�Wjr_r��E�qT�=ņ��|m3�#�B�����Z�Ô��gs)���k�K�-�������xӔ�%�U8EbZ<A����ɇ�� ��B[@��lX���V��V���$P��
��+"�'�:�p�9��B�Dt��u�[��;su}p���}e��-��Pj �
D��WDG�ͪp��[�����OWvĨ����>~DAK�v��qF�@6�2	iI����q� �9�_��5� ;0� O�E���+��l��'�ccӤ������=��A	%��dR���u����Ǌ��qK��'Imܞ��dR�,k@^������mY�S�p}ڥoG��8O�-<`e-����Y�����l]M�� �dd�77�����h|��X��I��f�R�
�U���O�4v�_.��g�M��{V+�~_a��C���� ��}�	w�_�Ylq�J�n�ȩT]@K� �H��L�P�1��6x���5-��
�;r_s}<��5>��*�Jm����?#r^��O�O�$�������	A��+e�@]_�ʚ����=�p�ELb��ԣk5�9��,�g�:����k>�bu�LB�ß�hx�Q*{�1��xJ����O1�����)=	�R�3z(�ʢ.B��5��铌^��݆�	�Õţtuq�n�00�?)#�Ğ��
o�Xh��b��ӯ�z�9de�?aPlR؋��N85]-��Zo�dẔ�����c��wj�Vx��h#D^?������^�.p�=Y��j���|G����d^`��H�d���W=[JU��?(�_YY�����R��m�m
��ϰҪʒ��U�.�z]p��6�U��29�D$��!�6��ΰ�B�ō����S��J�Y�\9�
���t4m죪�v2fۏ׻ѥti�����
}
�Fw�8Y�X}�����|+�RUhQ�A��6��Zz�EJ�1�����]0���^��>�����]�
!���G�U'[�����(+]����;fl@[K�L�{4�`�G"�� j��K�j��V0|0hB�|t��d] 48Ga6|����k��?-�X�r���J�x��ڄ�+dk�m�԰&���L��3�ݼ��kd�?bq��\�=��%_־������_@_�h�s�nȠ�����Ǵ$m�7n�����sQ�P��J�΢R�\L6
�Sr�<��I�,�몱/R�"&TGk`г��v)�i����zd7�W);Q����a�ۀ&�0��rLk��y�EO_�3���b��Lߍ�Q�n���u� wM2���Tf�F�&��dߎ�tfw�=�>8qv��Չi��i:�����i�-?��0�Kn�-�����g �\�|��V`2<��t�$��xgѺ�Pj!���E��#��:��Ț��5��Q\<�����pN���L$���C�
$���σW-�-�Xk�g�6:�&�m���`is96Z�W3�Ga�˯�\��4�������M���f�++�X5Ρ���'��g���?R+�c0��4ND�8N$�n��]�AӸ�]V�����9RvZ��M�tW�W��Q�	���,�N^���N��s�#���&��7��/2�Ⱥ��VEٴ��zd��% �w���^Fj}���_�]��z��`g��4�웗��?
G1��J
˺�9�=$��,��| ����P�gs+U�z�#4ֈ��<K�XP�gc��	�r >��|Ѕ❋�/6�*����	���Ör�!r��|�NF��h�D�4���C�@Q��T�^�#�'I9¬f�_��l,�|�5�*�|��'A ;��L����Q�����y�.Oq�+jC� ߢ�q�'��0�0�8�A^����1����!��[�/����V����s�dd	�[��M�omgcys������L5^өә��ݰ0m�;="(9&Iƭm̲�w����5�P4"Y����+�PTX�z7fE4'�9��d�IG���׵���=,U�2�L���m�d2L����u	�yq)ew�H�bؒ�٩j[|�E�LN^�0� ?:��[D|tS7��GO���K4��N�Q���L����B*z����}�3��A*�"��/9�W����FBM:�Z44 ������Ó��j�0v�hw��7Q(�WıS)���`�;�R02��� o+�_��צM"Un�2W���>��2ʥS�vs���oc=6%�p�l��伿��g��@0�����|Hս�uakm�G��\-�1żo+�<!2G��n�����"#�Pq�I�9wP�* ��)��Q�J'�d҈��/sӿ��e�3�,z�X�>����v5p�C�{_�Vc�7�:�2a;�CP�;����D�����y�判uk2)?k������.���j:�P��\��q|�>����ҙ��Ђ�R�����d�N$���P�+�b�@VTgκ� Ɛ�3���P�e���CE�M >Yi����*^���b��&��8�_�]M�_���w��*�n�Э]��up���?���S�
���zl�&Pq����V��ְ��	��q���7�z/�?�`�w@��g�I���Ȭ����QU��ő�R���v��*�&$}�f���}���X�-�p��{���"�=5���xw{ ��r�0{�;0�R�b �gNSD|8�+;w{M��0)̲8!Gλ�X ����5HvZՕ��'`�XR]"�&]�=9�!�� j�,b�=��n��U]�����7��[��ӯ[�>.\#=�K[(Bb�|)�����&y.Qz��:��q���
���x����[���������@`��pOƶ��Y���:.G`�Ā% 	�᭙��ť G�MH��Z�cc��d��E�v����0F`;=���!�� ��Vц�F/Ja�_���7��'c��?�J\T�$29lG�8����(��&k�p�n*B1��6b�2E-�V/�qDݘ��`0D�ˇ��``������ح�R�T���O'�6��?���X�o�#η鍢��{4 o���8 ��HO�3+���PзE���]t~����GĭJ�yP�m+���ܪy��C����~9��o,����A6�)\5(�@b��"��	���2/=%ڑ�\���~���R��;Y-��I��J�4,wR5�H���㼥�Z�zm���A�Le��U/u5[�_�oa����c��Js�d��̊?%:$=u1��N*�n��EW�:^	J�@��(*#�ޑ��o6��1YX�Z�a����"X��n�K�q�LS�&���u�j�\y��`�¾!פr���\�(�'���4f�/��Q��W�����;�,����l5����V����y}�k�ʦ�Rڶr2<�-:y�q�.d�"5�$���F��'��P���v+�5��{�}���o{���W�ުpʹ)�y"Y���In��T���J:��ya��M�ns3Y�b����Tꌛ����?ܥ
�	���r�7�>u�ť���1��v��T����r<xR]yS|_�;Xg�����3̜�?(*���i�,㥇� �L����e�o� �D�ї�`lm�k�+ԋ?\u�����n�ҹ/��DE��8>J�{�̱Ւ��[�Xl���NTw��.�����;�0���~z��I��w+�pn)�o7t�$�#�P��d��8Vh;���5VK�+�[�O��Z���Q��Ϟ�0E�ha����ȅ���u��$e�v,��U3W���殖��/9��������	�3߅�����'֛q�a�7�'nb8"0��z����曆 ��)�8*��,����O��X;@�ƫH�Y��|���b\T������J���j���Qœ�M��#ߖF��qƠ	S��VH`ae���܉���Mh�A��/a��=��މF��|�X��B_#r����n�B�P��
�:=���8]C[��:�a��)���UL��[	'��<�R�N\�V�<��7x��蔥�Dȁ��/�>����ނ7P,��l�E�Ɛ�<��9���t!�W�����;���F8u���Q�ї��/�Ϝ�����!;��W7$H[�Y�C�a�R�����;�K{��<��7�t~ןOy�0E�4&�P\���q�%CS�
Bk�R���.3��m�̧|���X�������Ɩ��Lf)��IM���.>Y^f�J��;�S�#8�[8�!7Ĕ�-K"��;1f0�7&��|�]�f�&m�ѹ����B�'i�P~�=-�}߇�F�\��"�?+ެ8�K���C��S|�[ᆧ�adUV�Gk���k��~�ۭ�XFi�ڂ��Rv!|Zp�QLb�yډbGs�Mtkr��I/}�/*$������T���J��7�͑Ҋ&+:$�-�hB���˽]�/D০��F�D�U��I"b)7mM�g�|�Y#�����l�x�M�}�(\�0���W)&L�0��ڜ���Ds{�.H��e��35��I�@���#�J���Žy�J5�	��1_��9	�â�7�����������7彥	�Gx����_펙Wj�ܰWv�O�> sn������U����ik�sh���C�������Ω� V2֟�*-�?1fDm�A�SJ����I�q�)-f���O4�1�|�$R�{Y� �]r�}�g�a1Vӈw���n8�������U{nz{��C��0%��Cr	����s�N'�K!���>�"35�$���^Y	 �Ї�%�E�cs��N]'����U4�@�ed�[h�<�G�nu��L�=��<�J�+�om>�_��i�J�u�o�5~��$�A���M�J�Ɗ)'?�)�R��y�H���L���
�ۓ�ʉ�f}䄌�}Y�g-�۪�_bc�(�e2-<���s�e�y�G���s����S����l"�U^܎��-�!�������'p����s%� o�%1�gC�ZN�$�c�ڼJ}J������OX�T�R��>�rh��N��D��ü`�r������1)�5J_&�"������i>�p�[]<����J{7,�*W�֤��?�s|��c�P�#��GHdp�9�F��I]�=3�ڶ�sBXi�go T���V�H��{i� �$�߶���5�������n�y�(Z�-��ωO^%K���B�A������	�Ig�Y|�f��ivcK���7��N?֩��J-pLj�@G�eC��f�y<+��(`Հa ��C��Ax����#J��A��V2�<b b-B<͉�}��层�6����O������E&�����|�͗����,��=�?r�@=�=7��n�yo��'&�(<Y��@�_�x��p�W�DZB���U���3��ߛ������/��\��z���(u@%C�d�� ����{�*�{_��c�(|Qz*�+smO�R.?�@�V�n,g!z��h���3�:�)����DŪ�7�����ݢ/�y�N��f�ƻ��Z>x����w���)�Yf�C�'*��^�Ϻ�,
8bhI�\\�d��<*}�"W���|�����f��㗑��\O�5�.5��"�+ΩW{Yߊ�+LPp�4<=�.%���rMHSRD�#h����P��N��C�!]�ުtK�BL#��)@:��h����.���A�����W�׮'�GU��&-:��6$�OD(3{����m�o�M�q�Dm�>{C���5Y�?�J��|\��/�d�Oȱ#��Y���ll��:K;d^�P:�.��r'i���C�nw����ŕ2�Z�Gܮ�s�G�Lׂb��F�����^�$+��q�Shգ�c�2xPi��]�F�z��X�OQJS�(�ˉzUK��Xvu�9banx��x[�IV6�+�^Pq�7�l�U��m�]Z%��Lh7��5} �uB\�k3����+4�}i���[)Uh~_�,^���U��=#��e�
C�kxR,S���/G�!ٻ��Œ��1s�j4���9�ܵ�5o��|��^�:�s��|=�[z� ��^m"~W3;jNi��@IȒj]��ʯF3s`��l��]��:�;�_��D֥��n�e�r��Y1����fn���Y��k~��?��c�hs��0��M5�w��@��1u��<P����W,���\����d�[ `7�O��b�Oh��|����T��K�Z�>tcâ)��(h��@o��S�3:f�W��GV�!��9]7)-D���߮Ə��j�����5K����g>�]\����n[I �(��Q�ߖ���Ɩ������@�5� ͋��@^v�M3#�xM��W���~���;�p�Ha�7�x?n	�踈�#��u���w�u鈋��i��d?��� _��_��0�>#,��O�)_�eA/g����������,�R)e�)o|� fr����UၜD�d7�G� ]����
�AY�w�:������y�GQ�\Ֆj(��� �;���J�>-�J�)�!,��TQ�5��$R���k��邥����Ws呥��M:�0Zۀ8{�ځh�R��	JwA���H�R7�ϧ�
�'���H�x����f�i$��/4���X��~��dȃ��C�s�ӧE���oH��+/�O��i9�z(�^r�}p@[4B�%-���M���s����0������A�Fc��I���F�?��!���179gI�C`[��)�^|��5�yLn�Ě9NV3v�	��㢛N
gA�ʑ��\����q�q��cCpQm�L��G2�	՛�H��۵ ��\H?��xE����vG4���+̬��ψ ���h�'V��I�Y�Oby�f>�g8��7e&���~�*�:�M ֛��«��m*��"qxriZ�Q,#.��@%����;J1^�,=�ܙ7�u �+9��Ͽ�I��%�@7Iw���R�"�R�wm�^��i��ZD�2G;����Զ��\KH{پ#�S֔�B-�l^Ǳ/��=N����_L����$9u'�@���i;�
�f�uݻ�%1��Oѕ�W��5���m���H;�6ƻ���Mk���B\X�w�7K�\��lҬ����53O��,�d\�e2�����R>0I�|����0U��R���vycG��]��L���ۤ��F�;��و\���� �{�2ٿ��x�7�����X6$%U��Aw�nx�8������6�h蝀�&����)_\�����W�L�p�s���,ó��y�q6�(�I�ʌ��`����<Śb �!OT��~�x�ԣNK��͊�|�<񳼎b�o]h��ئ���C �b���t1�[�-��c3��!^�r-4�;���Y(��CO�N!�V,qs�Dd�A��`��N�x�J�&U������g(�����H9��Y$�u�y�� ��������c}\K�\��S����?
waێ�6�E�H�N�Gu6��V����a5X�K%iN�vO�5����O�HC��r�e��!�UJ��ʵS3���Y��w���)�ЦVc�*p��NC b�f�`#���	U(��	����ذ������m��6C��}�YƏ=����6��E-�������`b�O�Yp�2�Q�H+M�Nj��k>]%@�`X�,����K p����ªcVI}��N� #l7��8,� ���n0�u�w���<�Y�$���������K��Տ�d�,�������;��Fd��n����{>��b����7��.D`�\��.u����������+�p�!9q�axl�(#����2�G�L����]������7,����cՎ����I�j��R��ؓ{�nP����k&Ğ�m�N���l�L��G~�Q�B���Ok^8f�+�p557.�?�e�9<��$���Ћgw���}]��F��p�i`�%w�G��9���o��G ��)�o�ӗ��>#����io\���7���F=ORh��!�8��5�� e�)�Ke����M�7��ʁ¡�B/���cq������7C���]�ԟ���(�牼+a����J �<genO�j�5�E�*J��O�lD;j���F���/�r��-(�	j5�%R��l�P!z�����,�S�EΤ���M�{�i�T���kuh���!UB��"Z�!7p��4��/�_s�XWf@��{ԫO"ˬ�ݽ��K��:n�q�x�Э#�i�Q�nNycStr�Cgɼ!�l�x�J���djh9�|� ��̝W��>j���<lN���)<(ne����$Zm��3��dԈ�������'��]���-�U�2�F�js���%�]|$]�'�S>�ܔ�2z��_bq��<"��)B�K�3퓉�h�kA\�ኝ2�"Jb�P�x��],i�&>O^�|�<A�*:t�ؕ������u��{^��ư���3Zwz<��oHDg3ŗ�
���֛�l�`T�ZT��r�Ґ�7�����~q�+}<�M�4�4��#�Hn��`�oɷ��ݠ$2�F��|�\��w/��Vͯ���I�/��k��%���+f8� �p+%��@���x��2z�N��dd�#���Wo85U��Wu�B���nn��\��U��v�������<���p�1��\W�+1�ǡ�)gq��h�Hu�U>��g�TH0`���C8�"�A������lcM���i�����*}�!���e�������HN7ҝe�`P~�g�y��~
U����50l�bgyT<$��o�4v�(1?�O�R�n��q�͋���D9� �>݈�Dva�E5��i��Δl:���m(��b��c���ŷ��LE���~[»�K+��������HPEw�5+�����5["�ih�����>gzL��"��&�W�\��,�%��z/�8�N��L��u�$ʘx{Z�ȓ�%�� R17^`�s;^��G�h����IM�ۓ��0d�DK�R19��K��ц�lM������&���hMDKΔ RS���+���$�e�b�h����.69�%���o5X�0#�:žnr_2Sa��Uק�k��z���"(�-/����� �=��u���q�ż\`�o�h͚tk�q}S���v�@�e5-�A}���
�5yޟ��$5�'H���Զ&\���W�8�k|��~�\�a~Mʥd䞸`N���~ފ;��zz)G�H��c�����N��mY<�Tq�9(��N��(!D�W[�U��� �9$��Y�>�ϖz�Qh)��wl��D�G�ɞHsH ���q�w/�u-�:� ְ�!i����9r�O��2bB�A��2�h���͡S���q��T���=$G��?;8�P�=�f�Gbjdn.ĺ1�F
#D��e5�&�1/U,�-g����>�hZ9_}����]��x��%�G�*ÜH�m�a�[��.��͇��#=��U�^HNT������`[�*^� ,�����*\t����{p���g����s�p_E8Dr�,����b8mr�� S�+=Z��u�4�����X��c ��-�f�6b���h�ɉ(�n��z�E	꿝��H�	 ��[Ϯ`�a�k ������C��GSGe��X���݌���+ϓ8�1pB*{]W��n\�W��×�8�=�aH"�%���I(�1���R���P�=��\�d�=ɵ��k�̬�GV�`vPD�$mp����Fι�������Gn�f�B9,�
��`E=+�;hhЛS�x�0z��P��*����k]f�׻-����ď�S˜jx�r.�}�M�{J,����=&��Z�_$��xs������+m��lSm%��W@��\�W��P���A�:�
�0� Z.������@�E)�k��_�h-�����.�iBL�h�5l��ě-\۔h��m�o����f}$%���-��
�s~��b�#6���3R��-�zo�c�.�g�=:-�"c�P�q�_
y�d�V����x��2��i��IC{$�E��,���'Ma�n�_��6���*�,T3T0�Q᧲&]��	!�e���`��� Ǔ��|��>�����o��`���_���28�FU���ΈD�r>�M�k����.��z��J��$�_���o�P�)x�BīLۭ.3��}�SZ��s�����}�9pܘ�6��YM������s]Cz��fg��FQM-��\n9!�m�R�_�^c�ɱ[�c?�P�c*V�s�4�:�7?͇�bƴ�ѐ@z~�<�w�q���t��8���('2�s\ӽGPP�&���	������	F�Į��Tn�������e3|Z�!N��O-^�g�.u`� ���療C��;��o�7�Z����?���k��v>c G	--���^6e�0��L��˾ص*�u2Z�ݠy�-ox;���49!������u��4*#��e�cݢ��Oj�!c'`
Y���U�4�H��8��;Q#�����V{r�_�E�WQ=�z��SYs�y�AQ���9k�e8�a�B�Bf��c�:� T_2��C7Y���pv�7� ��/?�`U��k(3R:�T�m��"^������}��*p�d&f����![1��ezb¹����*�zkm�i �8�?\�Z������R8B�|ł����的3�{�)��,��s��!Y��LRИ��[��#��� �J'����_�ߐQ7�k����̐��M��A(�F`�d�GQ[��!<���v�H�(��4�(f�О���Z���u�=��WAر��r��.h��(�p�E7����"�t���DJ����{�����x���l��r?�"���yO{�6�A��5N���r	N�5;t'1n����$@�~+d�nȣFpV�N;��$?l�����7�I�¿}���L�`��>�ٗQ�C��_?�Q�.DV�����G0K,��L886Ɓ�a/cIQX� j��U�ךv'Ӧ�U�\�Z-�{�p���� Ud[�o9��|��7L95Y�⋪�̳��ٌk�K�~k6=8��=�X!�l;���넊���/t�i��צ��B�'C��L�R��m�w�⯑3
gs���k����ᴿ���Dޛ���g�ę�h"*�z�<�<��VtM&����t�����27d���Qa��?��7�����}@���J��t��q2�y�L_gjY��#���x�㠬��p!�>�/S����wo?d	%��S�B���w?了m�f8���Dv.��o����΂u�f+�ywQ�����e�%����磟M�5q�`���v��Z\���m�s�c̦;(�f�M#!�W� ����uv:]ɣ%.ǭ dF��K�i�9��IĆ6�����h!6v']�y��_�p�5���NM�v�d�ZE�*D���'p	�m�*7ek��V��k��-M�׻��}����^:���ԡ�� R���K�����j+����:�S/�A�s��3HY��xy<\63L/�=6���;���{��0Db�$N�yb+�E����ȁ�Ta�
������d�̨��T����mQ�cw)\8�Fu�օx2F��c)k��_� ��94]�A�eb����Wz��	���]��-��D�?#�A6�1�r̔�a���K�h"���UӚ�;�W�\ʨ����N��Zt�o�[�`Zf�zi|�l+籎/�	�_����q)�|� ������)��(V_�Jel՜0�W#3���1l�(��)����d��	j۰B�d -���mQO����6��= ��&�侸�Y�}���X�Q�D_N`'d�����7F��;޳�s�b��n���91`Ձ{4}8O;��Y��o��y����l�3Z�(p%��*J.z �bpx�L��<��N���*
�}8��ÉM��b�����Lݖ�\'��2!�7^�q��5QZ+�]!���C��A�������v��UV�x�|�IHK�p��E�de�d�\�v�	�Շ����}XN��_��d%On�F1S��]r�%X>|����$dNX�ԡ<�\ӐáZ�6#	�?�KV�xU�k�G^*��?��\�r>�\	~#�6�_)e�<�eR[N6������SJ����^��G	�88��n,i{���0�x ������'�Z��MU��5�"t[H<)����P������8�'�G��u=��^�>�H�u�S��x�~����i��Fc̑�ƀ���:Ei���ۖ c�o�{dM�;ss��8���k�u(��g7��i2ai�R�<e�DϮB�G�����L�5���*���7��Xh\FV�z��Ҭe@;�v2��O�$������T�/��̔��Rbj)��Hӫ)9�z��
��F@"��Q3^�V���a���z�G	��������m �.�#)㯯J�I��;/�:J��6�#�_ �vS���O~�u�oX}�����4L�0�UC007+�Y���,w��F <���m�!�g/hPe6��3+����H��m
<��U�h��u������^�.��+D�ٺ��6�*S��F�z�z�{~H������qzg��y��`C[�~"�IZ�a���ϱ^Ȼ�����{%v�bI������~5��K�(E7u�w*��Q�����P�yy�}F(�t9+�� Z�-٨��xNƸ�D�c��T�v�c��$�#�T�Ӓ�(&�P�tp(���u�r�(Ii�>���2��c�����߷�
��h�	[!����6os%��X�<��f[������$����uQ��ּB�kC_2ݱ���h6�fwoA3�Hw.�u2�˂"��L�F���k��̳q,�!F!�lG!�O�kd������N#��Č��?�b7�Mhf_�3*XZ������O���9��b��f?�Ӗ���i�����9B��Y%(��|Т������
���R�+p�=R�SA�dj����k=5&;c��%Ь���Q������!@GY"%͟����F�__�8P쭞;N�s�;b{�V�����'+ˑ�'m\�x�n;�8�d�OJ�O�?$��f��=���8S��#�?��,�(% �T6�=Yѯ�dvA�P�yT�4��Ĭ��N�HSLZ����/�Y=�n�~�\�}%ͫe�2�Cr�avS봁(1��Q
��?��+Kd�%�Z����c}S�!�Z`��m`E�et�'Y�pxv��T�k�֓�!���F�@�]mr#��g�.
P��Eh}��0�+V
�:�s�aP�ܿ�I�Ć��<֨�L����l�Ỻ���W�Dp?҉�4Ny���MV=f��ϐͩ�v/?�9�)�F��4[�D[T�
*`�ԕD�(6ҕ3����l"A�Z��O�(�����(��3J���\�d��[���I�ϔ�_5�3�f��-�ъ�»t�K`�c��V�o''r��, �㡘��@��(~�����+�<��-�.C(��Ӆ��$M>}
�ê������y¢R���?�"�X�Azy=0�k��-Ҙ���NE�֒�z�)�%P�:���}� (��5���2{���$h:�85��t��g��k:��'�ݧӎy)9<�ѭ�f�
���D-e.��;���%ǘ����y���^��M7��-+�c�t
'�-��z��=?�&��G"]eÄ#��
��W@0��Ը���V��r�sM�������˘��j8C���7轤\��Ir=յ���k��2B�Q��5���#��֙3�����2K�ֆ��3�{��8������5��⮨�Dd�t���S꺰)���6=�1�K��a�$H>e�6�u�j���$���+���`�Jc��6�C�dD�cX�k�[/��uQ�e�g��}�˻ �)��AE�9i�����sg�E��� h �ǀt�7	>�N�c�%9ɏ�hZ7��Q��>��r��
{�Ȓ�|��@�"s��Vx2��YSv�3j�AA[�;�rb��:�k,�x,U�u!���mT���X�~�/�z8d?��9��_����<�8��U<�Qѻd�b�l����d�C�.��C�`��h9C������`��a�'2�G6���̂B���\���K�u��X]�0�y��*��tC�7�YK���7
b�?�g�Dݍeނ���=����	�Gn�G��#)4��40�©dk��+�����"\��$�_��o������n�C���x���O��	s�N��[>љ�B�j�D����^2�gr6�!]����٦�����0k]���� � �Z�ۄ�Q�� 'u��<�ތ;����={]�I�̏.{�:vl�[�,�<Ay��hL:{q����Ғ�70^U��Y \_y)�e��T��cH=�����X�8���N��c�|h{���_��^��񮚻�z����"C�x�|�	7��i�vs�u$h5�GF D{q����IEMR�"` �7GleiG\6{�����("M0P�" ���sPR{����ô,p���~�B8���E嶃�|H���?�]�j� R�I��y��Z����2�I)�@��8S�_ed�+��1�"���G�n ���P�O��آU��q"p_	���cV<e��j_8������\�-鬓[~�R��&Ց�)��y�]0ϲ�Y�K�5�.��;��V��H�Y�F��ڞ��Gw��F�g¡�v>���5���{���~a"�~C���o��W<A�Ɍ��p��/���{��EV�,B���Q�M	�d�6�n~Gh\>��F &5�0H��EQ��N�+#!���v�fU;8����'V�<���%�
~�{�,��]ST��X�T��B`a��G���1�/�4�v&�ud!����%tq��ٶ�Վ	!o���n�NBh��[��L^���e@oG^�����������Z�W���BL�ު�	X/ڊ�����[����FL��92���b&����jD�k�K)�OH�{ZFj�%�)�3ē����aS�����'"��R�#6<���H�<!ӛ��aoFk}�(ٽ���o�V���˱�o]�D
h�?��]$u�c���dt$�����Cj}Z�0�~���W6 Upkn��Ko
m���/��GC��gH��l����*�����b:�JxX�x�nc��l���P��8����gR�7�/�-�;H �%j�kZQ��+�"���i��@>Z-���l�R|+\͐+�0�_��ay�*�}�����Y/�D×������CL\��+���K	�]"�mE��b%�}P��53�ۭ�!�բ��+o����r��	H��d�9�����u_[D�R#=}��7�mc�U�IU&��z-<I��z�K�#�<�I;ԏ}M��V*ɹ�c��i��:̪�`���U?_�a�ra�>�g׃�I��I��'Z�i�#\��w�B�߲�!�M1� �TY�5���?<H$�ŕ� �Y��=�+л�phכ^Pyyۺ�e�ۚ(�5`OJ'��A�o��_,�bb8�W|
q�v�j�Y�����R<W�fC ���s:��s��/x����:�����hľSF��{��/�ꏯ�{�V^Y.V�-�8DbM��&�Άal�7~�W4�h�#Z��Z/M����5j!aO{?OA����㿝�'@(k�<c"k�W$w�g7�����M���r��������-ŘпɪE��BD4��*��11NvװI��5�߃�v��k���"p�-��uI�(��j�	�c30�R�P��B���o���-�D�+�<�0j=��,$���er�T`�q��Ь:b)5���"e@������½]9�/G��NW�z�F�AY�ٹf���i�4a_��#�$��k|�y��9��sm �>:<JZ�_P֊C�3pn��{Yt�5�`�@RmI�B�6�2o��%�ak�(���ʻ9*��{a6ǩ�M@"�P��T�d��,�6�X�uC��g5C[��r��]:�hS�a7��n��ռ�.O����B��T��}?hg�a'Џ���yw�N~sn�مwK���u��bi �HS@ܲXOKM��v���N�xv��ɴ�?v����"'���g2�:��3��Co����绩bW��Z�$�դy�6�e���|�]g�`���aKcS^�ɩ�Q���R�I�h�Q�C%W���AGY������m��y�; ��Z�K%~�D\����x��N�{o�b�c��-0˸�����3�T
4n�\M��̢�Fl����N�Gt�|�Һ�b��^����m�R0���3�R� ���B*�26!�ˋG�M�v$��/}`���X�	}b���N�~G�S���I�z��2X��	��AC�7�8��_���ZN�,���S���,-�$8�\��/��*��b�ƿ��M����p0���0>�.`'�����y���G)��ڠ�Km�	ߒy�ET�]� 6rH>�'o=�g��h�g�OD"���3�F R�Tv��Y���F�>-�}�:9���C���'%�m`�r����V�����y��@��|Ya�Ąl�x0����V�X6�%Ҙ���_��1�6����m�� �8� ԗb��s�^�R-�
��l����oYv/�5�D�Xc��B�O��ABPŕAHa��ɭ�~���@/�R�G3NI�Ib��A��JU��~d�5c-�i�w��i���uH1�}X�9iEh0�T�r��9�@KQt��]>��uF �1�9�J��~�uG��+�A���"����i��˦��!i$��ås``��u����WFr���u�p�BWS��(�[$Ki/�������?���D��O�dn2�i.(�#+4���6�E:��Q��h�/�vPp������Ƹ����:\ZXD���C���3ՌJنGTDc����7U��22�$&�K�4"���r0/�l�
і&��/�X�w�^ ��֬�ַV�e�%�)�)P�S�w�c���0�Q�ܬ+3���i���ء�ӣi�-��e�b��k�<󃖤�ς���^�˗��Mꦆ����5=IWJF(��h���@/���?1��u�T�u7�h|����҂��aK?$����yk�]y ��^.�N 1�RO���'b���y2(x���<4V���8P���TQ��?(ʇ�f�N��H����9O=��gzTv@�T�mj��&K"���L��O>����|��y��cY���(;�Cp��%��wϫ�	�7��|��n��X�\���%[�����[)�?����0��:�o�'�d�j���g��	%0d�Nf��4����r����t����3�\��W&o񎥇�h��Z�_%`d��&J��u���=�!E�D4hNA��Y�3��ś��/���\+�H���Y �R���ƐE_��6I^��H�-:X��=\,�X,������a���@̫X]]������Ad�B��������l�ʄ3�)~o���o7d�8�U���7��d5Y�)"��p,�4ߝ�¶`�o���"����/{Q�� wY\z���_�6�wt����)
���]��N���_�G�=�Q�D�o�5��-�s�rqc#���W�G���D�fMr#D�Aܪ����x|�$���q����j
@U5f-CB�PC�ΦN2"�J��N�����7�5[�v̟S��;R��=����\��9�R�'ص�3e_��1��$���eI���(u�}�ͤ��m�Y���U·7ع��q����/*%zq��[P�	�6	U�B��
+ȁ˧�6o�?2h53w(]�3�<-�;�s�[D�M�_#�&w��
��B�$�|�ƙ��K�p��T���1��[���	�4q�y-*���sĞ30/�$l��5]���)b�{s�GqpK�	�ߩ������Hh`Ǹ�{��tzB�^�*;�K�:�\���u&C&�sj�\�́E\��l��mH��7W�^."� �Ǻk�I���0�\�G�$��H �Z����jIoY����
h�:�U��x@���Z����P��
�X<*5x�X*�ErH�|���w[�Yp�T��0���E���j���Ć�ED���U�*)u�0O��	}�Q�VTm��֕=,@���
[�F��g���Lm\�k�<�'�`�(GJ�#��w�����|�TΈO�T�޻a���������ojy,B�q���=��P��\��QR qJ�H9��+jCdpsb_���.B�D�i����	�W	�8CN�ѣ�)9Se6l�$�L���/䛹�,{x���JpVyL92��N-�N����`��@l��~с������h����fs'�mu�;=lrڔ+W-�?1Q��_M�	}�^,K-3��Ayy����GI/R���	#�tV�hX���I�(��Ck�<%�y��t�,bh6��[v7\����~�zjt�56��*R94��hA���Zƌ�@�;�� ݋j�-�Xl��d�
���2\w%i���9��J��p��6��&�s~U��*�/^�z�h;6�rOb�`��e�{�:�~*�6D������P��&n�Z_�TW*ؤF]�!��Ð_VӒ���c
]���O�]���?*�i	_��ɥK�F՛ ��t>��d`I�S������8G�1Y�G��^6S�-yk��ق]��*K%��O5F�yM!�|�j�?�7���v�.�+�|z��!c��[�/�>�� $Y��.\�k��0n5\�%��EN�Q=!����/���:��Zc�
��
�R~a���P��EW���_H��:U�_eݥ���aV�>+v%���{���x��1���yRG'����_ͶSQ� �ퟸ�7p<���'2U��fO�4�-�f��ia�uĊ�� �������07%#��T>���!�O�R�T�³t-m�j�i����|7����K�t%���e
��{�Ly�) Е���B�	bo=fTy��o�1�DǏ�P�
�T��i��jq(.e�ֱ쩷�>�K����W��J���\���ݼ�d�l
�C�3$�6H���!�����l��0&
t����4�T'^��(��o֢�k
��1�����t=��yj��.�\����B�7I�-��r��uȌ�o��� '�Q�F��;JM�\����I:)A��
wRޫ:oϞI1��Dz;����#���M��>��(7��~��gw�4�	�*�<r����[���:H�*lV{j����O�-άe�D/	��bP��2Ka�I��!z݆A�V꼱!�h�=uo@�]`�>ȃOn�I�#�����V����!�}H�6;��e1(B�=ah)l:a@ ĳ��4p���ny�{ӢX�8����~���l����u��{����۰����g:Q���	��A���91ڢ�:D��_�~���!�o�R"����䗓A�Y,|��N���]ݪ-�kA�؟���5|r�o�� H(qI��x��z��*]��;����P`NA�G=�*�9Md���/�ȸ���t������)�}�G��a슏��Ҩ�d Y��&������0}�2�tQ���f$2c��չL�@��BE��>(˝��N,�h/y�W�T���� �%���j�D�4�^o�Q����J��N�D��J��/*8a����t� �|�gy�]��q���*C̮~��"����`������{"��.��O�^�42�}D��k��p��Z�w��Y��X(�wW��ndM�$��Z1��
�)p'U"����fAz�L7�wY�Se�h)=s�~�Ɉ��ܘrn�|e|�*r�u����J��6 �ӠEt��ט���7�9!�TK]{>���g�0s�?�������5 ��-����հ�7�h�`��f�|n����b��&�=����u���ݧ���Y�x��461V Ah�v����u H��K��D���k��g��L=+p����f�$'Lg�'�����}�#��k@�"���o*r�WЇ��+�^�����ɳ���X��,~G��4[b�*�1��ټ��Wr��K�hR�W���ٽlvy��&ػ!]�N�$������`�77u��l����.)tA���+(�E]�Ԭ�5P���?YQyI��לV0��'I�~�6ϙ�	JGi�(���N4
�-T3�zj�cj텶��m8���G���w���~1/�u*��N�Y ��
��%WX.Ǉ�J<��<�Q�~V� �*�6�����7N���Z_S{p|P�Q�N��F���s��E�/&�v�wJ��ca?hT�Ծ`�j�z����5�����S?��RrQ;�Й�0���1�e����,{]�>�skj~Ze����
}"l���߳��z���2�XXf�NA��T�_�0[8^pD�o-�x� �jhb�Zˈ�%��wq.��aԅ� �����Q?��>,.���K�K�5�d��x���`�~��V�Ӣ�X*����y	�R#��^��_p��wj����[��byO"��I�D�KH]fX����-�?9�ϧ��D��K���a�9�fnK�N1�Z��>,��b[���Ǹ������W���<�JuT0|�>$������@�Q]��h�DB-�	�j����ukif������i�]�~�2H	�ƙ`%Ɨ���ͬ'�.V�(�O�>!��Di:)~���0��(�ō+%��8�p	�.7ʹ�O�+6�ur�֜���yӾΆ"@�ƅ6 ���e��)a̓��6�/]�L/�����[D+�_��C6�|�C%Kw�xm�h	 ��>h�Ұ715d���-�q���3pwr!f��|������Y���[TnV=���_�~�Gw��E0�����Ė��N��eGS�2?w'&ʗ݁Zz�[�$7�����ܭ�Zl�&GuP�
��joƲ��d>K�P��ɾD�n��gw���	d�8y��j�Hu! �����}�M�Y�S��>}���r�|M˭x7�iAi+�yL��ǫP�(b�L"&3�1 �=����l�6���	�BS����Q�05��f�d��"-��T���|+ѹ�O�e�wiRU]cmi�n����Q{�;o�k�b/�CmIr���u����u�5Џ%�L	�;�Ϳ�8�|Pf,̝$1��}����������,.�F��S8�p���݃��������H>�Ҋ�xP��=�I�D��g�$�{�Az�c��`�*ܯ`Y�x����l�gG�
=&���\J��sG��'�+���|��eں�bN�N���!Z3�+`�~�%м��E���^��m3��� ө�>Epo��J�v>r���H���Ԓ�a�{�]{���:[��E؟����|�t-�y�GϤ�{���~���p��'���&5@�<SF`��a�%Nuhp��yH��.,
:���8�b�4i����9���PI����f],|a�u3���	�جA����dm���<���@��O���"
�ӥA![�G�w���)d9��3G���Q��dP`M�;��uw�|#.�I��b�OIU���?@�Z�Ԅ7"F�����vj�y�u�r����R�	�9L�,��:�d��q%����V:�~H�0����9��L��*�>���DڡZ�K�@Ğ��u��-x�h�a���"Ђ/-󤑫rď牢��8�L�!��pe&J0��g'�B�(�a�L��j�h�>��(9�\\�L|��9}P���(��Bp+�9%���j���
&n:����Un/�J,��y.�4�2�0GD��V3̎E�� �mlm��'r �]N��dabH%��X�:>g'B�	ltv.�U���c�Դb<f��_�p�%�A��Z݇Ke*�w^�{�|��Nr��:���`�g�AYo��/���xHSnqA�N�l����պ�t��u��\?�b*�2��xgC��H)��������2�l���8G������RRXC2N�ꯞO�#9�Z(!o~l�����H9���yS-Ʈ�⃫R@�7=3���pqK���*����]b� �x�H�fTp�
9J!�1�ҡ����1�}���e�E���$�pvU�MB������ 	rT�ʚ�FԂ�)[��]B�����R���3o�`�x�ُ�ܨ	�M�|��R��F���zQˡ~`N�Z�D8�{�BV:?�~� a�Q޲{��J��\X��z��Re���<�����ϣDw[�z˹�o�3 ���ƽ��˒��p���,Y��gY`k�{����6)��;g#Ԭ7��>)S\�'I6\6��T�9�AL���0���
�M��b��8�4�y ��~���q��,��`*�|Oą$܎�_w���a9�޼���9�T(�!��H�<+�A����ى� %���4^7Q��ɂ �Q�OlJ"�t�3�ٯ�)�l٠�CIHq��	6�P`���}�be���\��|${sߜ�ᡊ��%��z�~�&}�ȿ������s�C��%�R�s<����{����&�2}��yh��(u���>ߣ��@���3�ْW�Y�}�_$}Ogc����$�G둶\�!�vދ6���L>I�r5�W���3�ϯ�F�f��}�fJ_�<����Ԅ�Jx���N#�s8�6Q��v���%���@GӌG�8�ڸ�>��TωҌ�C�+�\|���H`�%'��M-·�!G2�a����3��*j�%��2!���Z��:V��F}��<�Ԍ�6N����|����z_>�\�R[��H��I�X��2�nT,rR!u��`i@�^����`N�,*Y��2��|V��	ѐNd�w��Y�T�e��Aǎ��j��9��pS�qs�
Ȃ��^K��CIt��3���(A��|KË~�������Qk�d6�f~�q��?�9F(K��'�,���~˫�,n�3���puf3/::.�;�V�jf�����#أ�|1Z�R�Lη�[�!����i��YU7��(��f�l�����8�X�Tyq,I(]�	�M���T᜙Gc��g������8���A�Ů���_���b�Y�#p��}7��]����G�,�1'-	*9��6̔g�i".�*/d|B]������&�b���1b����~`I9�N�ȝ'���'yτZ=�h��ڟ
SC@�vy�<�a�8�n�^��b�ѳ/�@�ۓ�B�Nצ������A���д�z���g�Y�HH�����j�C���n�ߟ����I�N�w���m8�8bD��%@�yD��q��%:��G�]J~!d�����>
���䐆¨<[vOn��RJ�v��!uB��@T�X�|���N��Z&��c���2_��P�)���Yƫ+\Ű�1梏��h$����K�]�Q��N-G�l:
R��{���}��"/�e�����4�s�_�H|ix7&LF�?�2�+k��E�6\��=׾H�t�#����sXgK�~�{��e����6���.���nZ>���������� fP���b4�H���f�F��s�o���=��7V.��q0�t�I�x|�X�ͨ=���K�
{]mE ��Z���Tג�k�h7��-��h��B��D��6����%G�yc�ݚP�L��C�6��N�:�Qo���;���{ �����;������iǞ h�;o��/Gf�Jg���$Oʩ���|��řY�_�u���2��������oIvT.��˗c��;�- �e�S'<�A��3zh�+�GN�K��uE��ᢝ�S º��D׀a%l�y^������r����1���7�a�x��/�7������.�����nȚ/��&�E'�೗����[�,�9�eh�ܝ��B�`�}��5�I�k���3Q�~�|�>^$�$���_����jͿ�V>�]��Qك���·�
��3�`���*�2,ڵq��Z��U�F������bEM�e�6$A�R�� D��Mˢ�+'e��#:Qr��j%"zp+Zx��l��[t�3f��7r��I(�6��ھ��<&��oOб��]��,��C2?r��11��=[���5���{��CC�s�g��Ǿ��ׯC5�;P�.
��c�5��ܙ�߫kMsb����mς3��#ڤ�*�Pk�#�Q��rӚэ�#�e]T�h��(~9¾�h�?-
�2k��Ԇ�P���zw�@�4bmnq ;���C�k�ʻ�$gؖ÷�r؈(:,�kl���y͗?T�9�2�_׵��L��{]�B��|Ȉ�X�Mm�x`$^R]\��n�&��k�����}0���	�����A;1���9�� �@��D��;d��/=����ס���A�	mmI��u�-�RRE�7-��V���R0Z����;)�rG�W.��|G�SU}¯ɞ���R��f�A|�]*�j+ɲH�7����]������I�xp�T��3V]{�-0�
5����]��M�Z]�_�.�����,蕛��]o*�ʷN/�D#C�D:��k��őM�8�_@��F9��O����;��&GY:P(�~��3*��z�`u���?a�� �Rcy���}��"<?�����>e�".i���0��8 &+��S��:��C�|�]ޚ�V�
ǃ�ԭ�@n�+�~8�G�V���$�n�!�ی�K�wG�uU����nh�g��}��G��&�RPlM?iz���d>��ܩp8���(><��4	,��J�[m�>��ݴ>u:?���5M�戴-�[x
����3Cժ�o��6�Isc�
j��/��qQ*$N]�l�����k��ʎ���c�����C�[-Y��&ܲ��1it�=����..��
.���V��Vp���-(�y��}T����!v1Ө���zʣs�L �	�XH=Vd}iƴ5������U]�7�
kz���Օ�l�z%�ȧ����X�]ƙ��| ?�l�qª���^�5��^��`������L�+���!����By� :!4]j�1��
?Ut�>�>5�����"�n�7�BoC�ƃ6��,�r���0�\v�E���R�q����m؀Zu�3�4�R�r��J(�R&�	]kq�gz�3^��E�B3�k0˭'k�m}�^�V������0Ҡ�w�z�5�N�L��V��TvL{�d��v�R �'k1�l�zҘ�\�~q.Y0�l�ɶQ���E�(��'�ƚn�H�N��<
h�TWt���G������Di��	����|c�;m���z��I�EP�%(��*����j��w��.}���N/�J�k"fu�yj�1�?�<����f�K�;`���';m���lܓ'�ċ/�B�K@�d�BG����c�&���N��R��s�������î�YC�~|���������B!��w�,�5?��f�=��8��¿
�5���h;�H�����iI�A�=�k�P��"k��MJ�I�zU�o���iT�k���9���
�D1�7z�S�s�{�s�� #�ʙܥ�ag��w�ƯS�f�*�u�V��`vO��m������V��+����M�j�.��$�_��_M��V�X����2"����R�U�w�)*M#{
��#aR�^ �a�y�ČH�"E��x8��&��]�2U\g*�����M���<�,�jM��f
"} ��볼ZZH����H}�k���Î������S<�I�ڎq��B��s""`I>,6�n�җ�6C4x�x�(�N`�K�E��*��NoOR�
X���ƃ�>�@}�d���Z �g���������������}��t��TrSw��9kr�E��[��	I5U�E�n��Ň�N��ɶĴ�{H+0�^
*%��0a5M��Q���j䜤�x��kPa��/6�T'}��jQ���˴�rc��S����wux_����RJI���i���������73"Q(�L�K�>�L�D)-a��&9n�x�?����:�L����O���Z��"	d�7��G�����T��ے��x<NtC�P��n��`��I7	�?`���Qco6���EBO"���\������㳬^����K��x�F��Z�`?i�9^~'� ��j�B�����j��
$'$�h/�j�U���/mq8>��������A����=ܠ��N���U0�����+"&��G'z"�{E�JJ)QL0���N&����@��d�)$Fgx' >��w>��'-ʴm�����0w��M�5��D��.�X�h?�°L"�X"�R�1H�Owf�K�	h����V��B �P�)Y��8n`5��#61��%~r"�:������v+6�+�Y�����˫*����0���_�1�Yg]���;�[�F��C;!ESo��:����6KHod�����<�y {0w�h��{�d��8t�nc�=ɓ�<u�^��q��A��Lp�O�Cޱ ��\�T���{�rv����j��q_q�� �D.CfP�6��>)Bԁ�X�}� ��k��ߪz
�B^�k� ��O��L�Xw�����E�o=�PX9�gV�a+��=t}�Y�1i{741�ڐ��g�bc.�(2(bgB���8Y�����0��o��jx	Y(�O�gC��U����e�:�K�֚��=Y����Xw���>�'!l��G:��<�txb�"�R��K��;��e-��`�~�,DZ�L`�RȘ��Pp=UN�
Ri9�29�&H2��&��"�~Iu�����8'$vm��}SF��ޜ ��
G8�&ҭ�W%`9D����1�<�}�NXb�9i�(X
;�!���]\�j�����Y	_�g< ����s��������Aq�@#��N��P�=���A��X��V�f�N�GI1P�R��SZ�ᦳ�T���QW�z�A�/!]a���dŔ��$���,��2u�u��_>��t�/��%wm>���:��>=6Z|vp	p7x�e�b^���w7���-��N�L%��}X�H*���dؚ&�V�dt�	٫0�P�(�\�EE��c��ֱI�X
L��O��/*�2��N�=(�S.8M`���?�U�o5��!y���{/���=�7�q/�fʋ"����*�7C :$mF��q�v/T�<Pq�3�Y�p�(�8Bٹ��4@@~�EV����+��Ǫ�Y�I�,��d��t��T>�qЮ+,�`"�"�⃖�����1h)�V�s��@~�6�fF��H&�wH�s��'�#"*%� ��H<��α/X�E�k�0n���KT�.�8�0�����sh@,?IcG�Y�S|��M�h��2o��E�R��t\0ٝy����Sc?I�u��cgnc�}��;���5p���0�5<�����f'	Uf�,�J.�v]�(��f��5��0D�pf��>[Њ:�o�T��O+;��I%|��׆<l����ԭ��P먜V��Z�U�Y���L�����t�̍���dc_-;��y�1R�ح8�)2gqr����jIB��������"��֐v�P��/����ˋ�r0F���e�]�"82���>2�^�w�ґ�pt'���wy���]ͯ>Ҳ�w��52*���1A��7L����Ӧj�. ����X���'Zw���V*֛�Å�[~���m��@Е��dӒ��[1���s�o)�á_!�FEzl��ʲ��s\�(#���H5�T��!B*\�,&jo�; -tg����íC��T�n���F��.*�XaD�K��w}`��j��ޜ�:���1��Wo�U��+}'n� �h�x�/��u�8.:���I������q�,�通]�g,D��ĳn�X��a%PWHL�%�Y����n��ٗ^B�jS�K0sd���d90lv"�κ7!�1�$���C��g�pP+?��.����E>'�R�`yw�6$�ZdK7�Cc����~݆�	�/�����%-�����+N��ꞈl �na���6����-b��2b�gNA W�<Yx ���	Pܩ�6ٽ$Oŵe�ц�ٚ_B ���Y���2.���>��n8]K�$�"�PL%��^kt��C h���_�<ߐ�E����`\
+�^�W�&b�A�>1�����r�{+F&0����T>�sƸ/j�7�����>���o�~^V ��}��u�'I��A� �ڏ�'i�����ˡ#��wzZ�o�e����AwJ��I�  ��0V�=..-��^t�����܊4.h�1F}�����W^�J��vK3Ҏ2���_'f�mX���KH�߹�l3mO�у,D����{���F��<�oYU�ZG�����������K�Azڮj���.\tN��^0��<b��)w;��B�'�9|4�l����6�"i�����8p!���gg�ʎ�p��n�V[ˈn�����N��y."_�uţw�/+n4���ݛ6�`(�$?a�!���C�Ǫ�qn�*���L��8+G�����߾�T,͏&?ұo�r�!Irb/�o3U�_
e�y2��� "��K��}�T�su,�lzp�ͣ���h 9悘�[M�B��H�����
��W���O�憫�3��������sE��i4Ҳ��|�'巉�hΛBܑ��	d.O��Ț�dɒ�g� x���2��pv~�ĝq��"���D�U�T	ŲPYѢ��f92z�T˺�����y�)a�	YVO��z��.�����_حP�o�D�zO{L�y�;��S7z}j�����ξÇ���L0�N(�^�jV�?k,�T�M���9ا���>��S��e���b\W��Ӹ��q�O͔Nq�����͈7�)���w�Sd���~0����T��jd�xh�3��o�-��8�]	%�?�+[��]��ݡqR�D�n�ֵ�AY�8Ž�v�]��#?��e�A>" ��OJA�!�'���o��uך#º���~���P�#�W���ޘ��m��U�UȻ��c�f�g���7}	�6ĳ����_�� �l�	LD���s�w�(�`�U�W�c?�g:�d�G��\��=������k��L����R�Vo�Wi����%���Tq5��{i���C2|b��灅Q.�G�N�_	�����%69�ZޞX�s���^dҘSs�A��k���'E��v?�Cq��U�a�C��]z[-��Z��s_C���a|�*�v������������%�V�C�����&@e9&B�>~�=�,���
ADU��<��K[�5RrL�n��x��K'�}�!=�S��O� ��;�5[;�I{n&�����n�+H��[����5j�
�,5����g�e�C���˾���iST��@Q�{���GD�
x� ׶eN��Q"7u��KQ��3�B��4kM6�®�_�d�)%B����BoF&+��1�D�Pxfe��'��pU����3}v�Q�\��3w��Ym?0oȦ�m��h�wW��ͤ���܄����)��N�ۀaQg�E��F�XbJ}g1g5�����n}���bˣ����h��ޞR���~l��Vx�ɫG�h�&� �VN&�s+kc?Բ��_4�n�m�Վ�D�P�]�������h�:
����Q�[���!�J��-���'W-uǄ��r�fOPT;ag�!�Y��	 ���Q��q�4Z�&C��g����<�Z�r��)M�9d�s�e%��$��>�����T+�����
�ޅa5J�ރN����"��Uw�^ђ*geB������;w��C��Z�T�	,�tZg�T���bHF�5�E�_yӵ�ʄ��_�������Ț�z;�Z�b�1&"UD�lϲ3�0.ے��#��?�3&x�S�puXߴ"�{2o�m��@jZ�6n*��q�SV)��uj�k*Xyh���*�|j=����RU��.	E�h.�cz�^K5���F�J�c�n������J.}�<
���<��XE�U\Ҽ�IRX(�%O:���.(�6���v1rU+ �`��@`z-�Gh�_TE,Y��_w��ׂi`b��s�*�FP�\JNr��):�`*�JD����%A����k�Hz{�뚭%�Q�*587y������MF�1���)[L�/����]8�K?�/�~c� ��;�.`�A��ht�&(�n�}�8���I��_9c�9P���b�k�;0�TF6�qF�3 S�ൂ5��X�&IEБԛ���o2�:��,�a���Gz�8�}L��9��,ZٟR|�xU��Ո�����uAr箈Q�Kϊ?' 3�p6�zx[��X�_���pL�p���~
YG��j�lm�My�ϚU����$�d�&�X��A��Ӻ�����h�ɲ
 yH��	���R@��47���`�E/7,��������P�[�׭*ɻ���v������x���x�^E=�vZ-��2u����x,.�cq��6�t!�"{	�X�+�3'�d�������A��Ԯ!�YG�Io{[�D�gsZ㳵u�-�:h�!Z��(�UC�0ȏT�(�u=��q��g۪A%�#;��u�����joJ�����,c -ug�9@��zt/��N��BD� ���/T����/���n�8 �v���N*��_g�k'CВ4}�_]zRs�[gT�b�C�J��1O�H���[��6Kc�6�]�̇��]$?��ֳ/���D�^�}j�P�h��������m"�6~����*%�i����_}u�+tg܌	B��@9K��G���h�YP|�j����s�4��o�j�5�[)�f���Y3}3Ҁ�/�nq}Că�/���	��J��+,�t޿��$
���,��wyd"6�[�"
��Z�H�Ve�Hָn�7ȸ�Tk�V �pk�+f��~HA�����=���֪%����ʒ]���'bÃ�yw���VV'�?ݍ�>�j���:�ݐ�46��Ń�"������#��X�Ŧ��6��"S�<v��i9�K�ï�,��h�h^�f����q	�Rd��7�N���ԙw�J�_ѫ���߾x�#��$Ӊ�p6���]�c���>H�Xp�:���s����{A���K�N,A������3߁6��o4���,��S�R|1��N�H�:.��F<\��<Yjқ�ʬ��N�*����p�*`�Y��$��(9�ߓ�:���8I4W;Ɂ^(}���O��)w�;�� +vi���y�h���!��e�i�L��Zrj�4��;�?�]Ԓ87O�D�t��k%��s����۳�u�mp��c�*�R�WQH3��ؒ��[m��t��RH´r��5�ڦؤ�F�Xl�UUkA3����%���-~p�����
L�\0wY/�d�4v����ah������ѩ�9V>�4P,szӚK�q��&4&�`���%�R��1��f�cĝ2%#C���S��7#[+VM>zf���j3�-5��a����rE����|73~[��)�6t��zF��{`�{�dҕǴ�SV�%:r�=�s"�܍kXs�.	����7���d�݈�#�y^<���߼�c�	K)���x޲�To���_bW�ޚ�>9��P���C�� sU��'�r��h�>Ԇ�V�̣� ��nYjh��B�%�����ͧ���We��<p�thGݛ]7;\X�l���0���Ǭ�1`8ٷ%§��X�j���
V�e��N��� �ԙ�����M�>��H�k@Hm��+��M�[<��c��B�6����Q8�^I0h����H�{5�w�b��yگ�0��%P7Y��[����n�h�0G� xrem�����8_X�5�W�+��=h�����AW���s�=�	�q��!wC�����B�&��X��h����bE/�����}��<ͼ��[t���ڗ���cb�=&� ���H��G�vռ���`��@ٱy�����F0|��B �_��^�~I���:j�UkN`�*�Rӏ�8O��vr�h�k��]�`l	���V�b`}�&��I0q��6��g��d�L�lڬ���[���y�!�A13y�HXfW�K����@?�hࡵ�L��9pr�g]/w၌d�����&G���\a�+��ccr+ �<��8W�`w|�N@�����h�xy<(��r��^�(��?�#G�6*ZQ��c��B7�
F���XY_���R0��m�F�a�������2;�V=���`}���Hb�EJ]��!����K [?0D�]P6�h"���ƌ����E��|�SU<�rW��@����u3^�dN�� |C%,��^���H��xe�_٪( ��ĵ!�����׀��q���)y����3c��\�j%o��gJl��R�[�y��>�8�Z|sR��:N\�ڐsz�}H�)�K�c7l՛���m$�Y=�/_�.�=�IFwc�i���bp#pG-� k�c`��
 ��D�������!1��,� (���5�[a}G"��l�R8�����nT8��:�q��*�����K2�,Mń	�y�-v5X�k��-p�� ��ouA�g4��ߟ�@_h��v5M�H����
���!��S�	b~&sGn-}m�����
��k0Sor�{��.�d�=Ud��I���!��9�2�x�2��ϗ?�B����>M��#Q�6U��ЊIo�J��0���%��I�D5�'c�p61GǓ�ULh�3G?u�b����cC�@(YB������8:ɴ%K�wE�
�E ^�8�NU��/���K�s��T��n��鋪 �݌�W���v:4O��D�<���}ճ)�{�m�JG�������~e|T����*Y�u�+xm 5,-�gR=\�/אrXCI�'h=���Y�\���dG��@�B}�T�!��i���>�-��ڵ���p��(.���VM�h�v��>����z*��h�j�j�f����g�T�{�:p
��'����1l����7���jFd�,2�N��<L��;��-�q�w(K�>�T'��W_R���G��q�!���{>�]q)1����Y�@������B�����^� �|J�a�/��ថ��T4�5����kxGiz���qd�y���)�Y��R�����+�9"��_ܥDR���?�{wj�����������$�9��
���e>���C��E_�E�Ԋ�zBJ�>i�c��|R��a���^���݊�$hʦLDB�LBi�w�d���wpo"W-6���2-����To.v�p�y����6`���!��}�T%	��G��x��	���'�j����}�>=��G����И�t�EH{���;�ѐ�eW{B�S�0g ���uU������C��)�j�FI���Q���/�y�XfI�. Z���>�(dh�#H�s'�lJ��+��s�>�-D
��8�O��
	Z�Q��q�)0�{�a�y?A�W��:�f�H$V�n���N�Jc۵�.��;�CA�8��h2�Xz+��ʐ��ٳ���~�b!��0�?�
~��	Δ��VT�;�{08AŬ�+��Ƶږc����1����z���ݙ���z��yj�!�3��3��-�o��Q��?���,^yl��>��Ū>��#�]�{X���r�_!�Zy�.�����6���:�;��%��uo��0�@�Aj�	`\1V����^��y����%��&z;�О�i(^�x��$��X㉼�����  ��k���/b[��j;�ĤMj��>��Ad�ad��貫)F�Ϻ9����U�(�W'�M�4�0X�=��E��j�؍�U�/�a��Ʌ\�M�� ]i�uH�f��kqb����g�F���!t'ڒr�n�4h)ۦ[S�ᶩ��ԅ��L�&÷�R�mU��0�/(a�����>���5����iRW����s�@��3ȍ�b e���SΪ&�#�t{�$�uA��u���������I��8)w�	F��_�J��M	R�NvF�HTx��z���:X�g}k���G�xeJ2l��TN2	���j�~�X��N���9OP��9��]�F���K��}yk�ka�����#����߼��"�F��~v�E�;�"�'��4�$d�0��Q�Ј��	WZ�}�ǯ�P��Ւl ��>�L��\�I�w�L.�y��.�����t�H�gL��:�dz3Á�Ro�t��'U��dю�z�m#�V�^k�LO]5�&��� �ǹ�e���c"�YW��
ǦWU���XQ�� ���)��<3�Du��W���e���?',�nŤ�ڸsE{�SsaA�(���g� �l�*j�$c#
�q����.Az^�d�b�E��[!�ɢ
����]�n*�;��C�
f�v6�R����5���kS�����EV��+�����H&�A�1�W6q٨?���>��VdC}ȧ,0��"]E����!��k�)Of�S�#�Y��D���)���$2f��"����m���	hI*<W�{r����������i�z����#t�}�����;�78q0�%��U���Wy�?V���῁c<�rP]��Rc�w���V3aF��WW�%���uI����LqO:���87/���d:�'��kI8.�" `��7���T^g4>)-�=��2���2������<�	��_Z?�6�|cXZ��D�W@%��B��,���׿�
�|����wC�6ԯ�\}�b�61�/
�HB�G�|B�8X�LM�GY-Ne���-�[��z���1)�*�
�T'/�
uH���T��Z
�ϸ��F*�����)����;R 	���Ǩ���L/��- �������X~������u���աV_#T�>��ȵ��MC��;ph�lw��D��w%��1{�Z�M�u-�{#�ve"s�Z���M�ɪG��=
��m��B%�5G�q�ͤ_�nj�&R�|�k X>;�t�����{UIa�"�:jH��8�����:ve�"X��՝��''����o:ɖL�4vY���A�kG<)O���Pr�u�y�D}�����Q�ɮ�?s���{�SguE�'�C�hl���=���6�3��6���ˀ�0�_B,��K���J�/˟
����0ܼ���rc��7YM��9����!�R�����&n檷7i�\��qz��N�A���L�
x\~���i��o
�<*�Q+�u"KF�n,_��EM�MQ럇,�}���!������C�6?����NI0 ���ke[�߯'I/}觷�ȁi�OT �,�#ih���)�*�W��wݼM�_w��N"��p%OWB��%9$������)uڿ9�a�ѽs�0o(�h���gR���I��I�4����m;�`�q?�ب���]�M6��=DI<]E�Jwf��O$-��zy+�Or"������f�iUTSx*���o�[��%�:UɁ���tS�m� 	1�ڹ�>��M^U3o�5O�##?���*���
�����h��va��`OUYD���A6D�圆�"��d�ƕR���`!7Ei��d�0W�fK*��B��z�8e^!�2��	O-�+\�9��\^Iݗ.�A��S��iT���e�}A��� �;Ř�����w�3'�7���.�j���sJ�U(#�	��e�jR\s�հ 9C[Ê�����(Y�X[� �N��ʏСPk�a����6D?��3���r���>^2����R�l�XJ����`D�.��F.n� =���uy�A��wr����-�7_'��j�E��]�S�H��:��{+T�[����>X�����f^�8c���!�y%*�v�oV��G�96z3���U�'Y@�5 `lՅ{����Cy��m�0��'s�}$��9��
��[��|�� ky��M�I?gē���}���5��Uj��1@�Rv�5D�O4��|�4nף�̸m��2�K�c�ؘ�Le�@ԅ�jtԍf��/2�<�	ܖ�*(S8���#�"+��"��L��UM^�[��0(S��yT�x^���ý7��ߘ�m�ʃ;�b�����eM�H�i��w��/��Ó�ub�Ѳ��c�;G�왛�(�851�/)R�������z�����{�����K��tf���tl~[�[���X�#
�ņd�W6�� ԧB���WJOd�`d\G�2sc�<ۯ������/k�\L�2R)�h��Z�� bycK�!*
2XU�<�7Sg1�9�3�jE��9w�D��+�u\�< � ��S�|ɹ�����7P�a��<>���Mmg�fG����De
0��`�Y=�XTDS8;�Ӛ'e�r�YF�oE����3�ʹ��=r{�Jx�����5�'���DY�XY�cw�;����&���^������̷e�ޢe�Y�+�]L�4���_��cض}�"���k~�� ����J��i]�����㛨�;�Uh�yC�)��d�ʖ�P�W����)�O!GZ�yw�<?������N�.�B��ÕDa.�D�,��QOb�E{_K�� s�p��e����~�v?�����`7���;���S_��!;���x߁]O�����"��l��nr�r9m�?��YJ�����f�`��Ƀ�������, � G]ev]($E�ñ���$�c\y���F��,������:����f<��~u���?��E����+ek�4��,(��* `#���<�~��c$�O��c���q#x(��%_O��!�]ߑ����|�m�v�!�sJi.��Z�����iY�bS2��3��r����_׻�?MvˠA"+�=�ϣ���$vVX`�f���^(lH�e�`M�$�>�"ن� R��F{��-�1祎D{�&��[aJ�������*������5/��`�K����*6�`t;r��!���=n��*qʳ���pyt�q�����4�&�������;[��*���,"����H��0
F��k�/k ���u�CZz"
g*���?����O�n�E ��[A�w���z� 67����� �X���Z�-�,�hA%eM�`&P�>��JN�[Cx+=��Wii>�����b��D$�t�3�����ÿ{�1)PW|[�{���m��d��'ݍL覀y(LATS��@Gq�(�E�?�������\�>�Z;�H,�~6��8j/}�IyrQ��^s����r٫&!�Ő��wBԎ~�9�Jp�'���6��ھ |E�D@�!�2^Z�uJ ���[�y:��v�B�%y����4��	R�:Ќ-y�Kh�}y%��T�Q����ԆǓ�B2k(N��լ�Ū��� ?��鍑�u{�F�,F��!����a�5c�i�khENY瀎��H"d\d�,�(��W����z�{U{y��&���¶3��w����ND[�'M\�ގ1'Ƶ�nN���x`	q�0�<uK\�q����FđbW+�K�d�{���ݝ��pk5���?����-����-_�J��u��*�wE��T����,j������I�)c&ʧ�-A�ů�j���o��4M�hF�g�}a%-�/�x�0BN��$�*_�Z��aB�\Pv�k��P=��r�B�E\�f���b(�2U��5Jt���b��ʣ���Я��8��]��z��G���� >�N�pAw�G�k��k�Z�JXF���(T*��[ԇH�1�<4Q+�?<�mS�����޲�0��X}�KX��ꂔk�M 4FD��V��i�O-��`��[�Q��7%#Z���>���d��8�������,M�
����xzv�9�SbXOݓo��Q��s{w��$O�2/���$/�3�1^��>������)DB��P#�x�%c�ٗ��%wJ���B.�c��XN�kM}�d���n6��h��5)�H$¦����;ҝ9���pH��������T%q��� 62���2�������W���%��s
�/}��W�tPm�����W����N�\6�p0BFm�Z3��ՆӚ]�/`u��;S����/A��"�ZUn�����6}ll���˾������fh����9;XH�t����Iu�o���+�����5-�\wp�w_���������3��E*B:�2��?�x���Z�KWgp�O�bxJ�W�'p�%��l<�Γ�ut�<��-n�Y�yE>)~A�x�A/�ܐ�Ո:}�(��B� �0Q�e	����>�~�U#f0V�G=��H��7��~oRc��K���uH��[mU���m���@5wB��qR�9��6��%ִ�A�n�(:K�vZq�N�J��z�qX"���H T}L/vB��%&�Ԙ��$�{T��������I��eu �Ŗ��pE��-�i�E�br�ze%u�~7�5���9�E�^-�/�οHY�VУ� �vTLv]�cJ�Me�X�1���f�W����M�:����ʹ�}@�0�������Pq0U=��HK����}����;8��}�(��t�ؐ"}By�0�iǾB�)$���^��QO��~;E�wS���MmRA�('G-�����P��M����=��;�S����j�,v>�z�8�Hu_ܤ�����;��5�X�yf��@�Rs�EO�����vA$u0xG=5��m����ۼ$]�Y���E���-E?���*����~�f���.�#�|&��5T��à|D}wI��"k^O�p�[��J'a��M�v3P�d�z�ZV�s�������|jh�ߙ�P�Q�^����AGMr�6�q� 4�^��-_B
f=9��@���F��/#�Q�m��"��+��UEq��13X����
������m;�Y�BK�JYt�iv��[x�����G�%+�1��r2����i��*�Fh�Ԁ���x�D,a`%�<똗����^Rǂ��%XI%kٴ��iZ,�~�ҽ����\SD0v�ʍ79S���O���0_�)]EN�P*��K���C����+2�~���3�q�Ne�%t�L�x�g'��%�Kw����_4����ߞ���q/������*�+Q���P[��长p�<烕X]f?׃�ե0�p4�6���d��?����S�"X{���Y�.=(�8�h��ru?ejm�0��ʃa(xW�����Z���J�G���f����{�]r�^�%^Ev�Zc��-�	�D�}X��4�9���M��p�ة��\�Ï!�:v�Ը��X��n�d@�}k���T}k�mg1�bY^�@��a���xe3+�OFs����eC�SW���a��y����{�x�]�@3*��
}\i�%]U�5v�d�۵�+V�����JZ��M;�ӡ!��_M�3hT۷��@���QO@�1�r�4-C���R]��"��A�z�o�P���v6?m ĄF蹨�/[1><0jI&�@�hM8_�n��{>�9���I4����Ю�c+�����
�
�x��ges
-=_��.�G��9N� =7�s��Da��@ΐ荀� ��"��3>�q���r/eS��{�d�*�O��/ƀg{Y��`&�S#i{��j�6�#��A[R��ϊo VA��^:�e1ᐩCP��lO U���O��J�~;�𧇌�[BR?�����l��	�R��rţ5��1���3�@N�<�F��]�	:�x	�>k�1ǎlk�c��y�Ӥ�Z��d�?o&!bM���?��w�K��>z� 9�`$',�üxH�X�ޫ�{,i�-��R����"��Q���>�DD=�gc�`���e���"�X]/���ӷL�L��U���?k�el�}���V\_��.��3�����Yo�_H݊/��ݍl��0��&�'�˖'�=�Xr*N�k���#+R)@�2FG�*e��J��y���j��Sc~�C�W-)6%�5������A^4�lE�m�_/�B�)�zYLְ<_���`,�r��#:�|�'N,[j����i�K��#��{��Ү�������V�|�.��+����
CC�茅�=X�i��������]h��Vv��D)�x46��3�^eC�t5j�P�r���̳ٻUT�O ��M��j�DG�hd?�:��cX޷�T�\��x�aj0q�9�K�,G<���s���ںh�Q�'�_�]���t�l���r��/o������E����*lQU��yfa���y��ݾJs��Zͻ��^^N{qlŖ%��2����C�y1��}�w׈�쩟e|������V�
ۯ�۫[�5|E�],�|�Z�|�)���s{�0�����W�r����EƜB���s{m&>��KN�Zz�OG����"β��a�A�(�csoV1 �(�a������+�m�Ή�s��ɗЫ"�cߝBRʡL���5lio��A�Ў��h���LD����o�W��4�-�YEI7�����%�C�5�M�Գv�����W�1�}X�ט(�q�)�6�x)���_��_��&�5�H�Ǣ�4�ձ������'����)�+�&E�UE/c��\�w_�t �?� A/�M��&��Bc?Yu��$�8�"]����qt{-�����8f��,F-%�ɥ}3`~�u��y\%lUK�
��[�Ee�W�׺3����v�,�
�Ρ�a�)�tqep�KGj�wZm��[5�1�ʿu�Y��!�2J���F	�\�m̐U{���+{?6�
��Y��8;K���S�����g?�]��鴸���A�(7GJ�x%�;���c���O;�V�⎷��Z�[����G���œ(aMr�Gh�	�r�Z���V�x�8\iU{�u�A���Z�FJQ��➏4-mF��SYqE�ķ�X�|CΚ�8�45Qޘ�g��%>p�)H7�1�龯�=�v�}�g�RE+Ə��E�J-�����g�rW�bS�EALe�����v���NU]��o��A��QL��,>��u �vc�q[6e��z��'PjjmW�sS	�#E�;�f������|�TV
��^��ǎ}����<�"r#�B��Ѭ��<,|}TȮC��i¦i$�� ?��a�^�7G�8���V<z|��!��qJº�-��	��`Ʈ���F�D��n�r�4비H���O����D�q�B	7��!��1س����F:��G�'��eW��% �vvZ�fG��5����Sl��_�J/�0�7�,F1�Q=4��;ʑ��Q�P3�d{
���RX�MkKoqf ��10`��@q�D8���AKjpGT�3!��o,g�&��Q&޿Ą�a��oJKPNXߝx��l�Zy>�Q�
�4{w�i)�培v��9�y��ي��R�s�O�������z�fԇ4�>�K���6�ا�M���Q]����5ʾSͻ� ��8�=!x��N��%�.q O�@�<�_F��.B-'������%O�wN3\o�ˤa�j�#t��{�X3E��Ny�G!��<�+����3%k�_&A��)K�i��K��/�0^�&�\~3��WH{:G����w��7��:b���=<�ߥç#����x�	~��t,�J��B�E�P��6f���S��aL�홂���{d�Ac@
R�;;_9�p{Ƴ���|8y�:e`(�h�l���>�O�����e�@�ַ�s�q7�*��6z�b?ce�H�aÒLn��.3�Z��U�F�,Qq�}6����$�t���~� b��"�����*<��s��\�)K;�i{�`8���lWxz����JM䔭%"5H�l3Lgj��g[/Ũ۞�׮��{ޑY&�4s�.����Nu�ֆa�T'���a�������Dh�u~Pq0A�y~�zÕc���w��n>��˜��ܬ[��obhV �q+ �{�W���;n%銀gi���۰}Q�`Ӽ��ڗ��]^�qn���Z�)���_�6/�,�ƢW�8��N��p�6�W���w�-���]�g_)�y5bΊ߾���޼��3&�� T�$�Y7�F�U�	> ����VT�i:���܉8�gr��nJz�;����B�z�Iͦ�e����)߆~nd	��+J��h��8���\���q�c���+��`��o��⍽l��Hޕ��Bΐ|��X?��)��-�w�Y����T#�䂋F�T�qB3,��xRw����?���Mi�������߹nR�*�a 1����qC-0I�=%;ι,���թn�.bdhC�0W�o����R&��(�Λ���9�ZQY,
;G٘��?��oZ�.�t�T�h
�m5�j�9�Qı� s�T���Ø>����HƁɝ� ~�O�cd��"�T������}�^4������v��]ɜ��Q=�8���|!��񪣫 �'ĝ!6���k�����5�߇�@��Î	��VE�%7�^��GF�^����X�<�"Q}E�^nGo�q�^WX8d䕓rEyR�2��]Pa�r�s����j��Y3���<�:�Ԝ��,w,;���O6tŐʹ���2Y����7N,�V�o��R(:�H#!� ��m��\���i
aݧO��������Zإ�ٶeP������X�����cӼM���͕����1�B��	�]D��<�k%�<#��.'}��d�uw��ҏZ��K���s� 3��<,���4�/�!�B�3�-w>���I��q���b���̏�p��=*��1���"�y�R���
Sa�i$���S�vQl�z��D�C2�j�"V���5��&pq��2����x�$}qҰ�W��	�Z�(��Gc�2�Fð3i��ڸ��G>�m�~`Ȋc��ޙj(�������1��c!lG�F�70n����c��<@*{ǭJ@�v��X��zC/��5����7Ǒ�Ν�������*8��EO0&KZҡ��2Uv�� {N�X�^FP�E(.&�2o�z��:_JP<��ff}�t�5�z�WG�+gA�*}���Hm�ƹ4ds��~�c���=oz)����r(�qΎ}����.��}L�K��bl�Z����$:�~��\p5���ӌ��%�����-u��,�2_ C	���ƕl���6��E�V?r��H���S0
!B��j��ixeH��I:�2
⛻K����X��(�y�8C�m�d�3%��>�����8S;J����W��+�v��jW��@D�α�N���r�!&W���n�"޽Q]�1�,WVR���Զ=J0�|8Ӛ��|"	�|�ߊ�8e���ГO�Ō�k�	Ig�3�jY,� �j&���/32R�����3�	�L_���� L��S��Dǜ�V���ږ2�-��� �$Wb����������Vc���Z�Dیg��(��A\�#���ϴ}6���+"����9��3cάKEx٪>�g�-%�5���PO^�H@{j�jSf>*�|�d���'9*�,��q�{0��d�X��ͅ�?���4iv[Z�ː<�*I� ���>j�c��<�!�~hW�o��"o�S��@{�)��3^��,�,,�4�c�Q�ۘ"�����h�J�����璾�ev��?�/��L2���[Y+�|��
�!���.}j��b�q*{;��9\I�#����-�ɶ&��}�:�j�S�>����*[Q7(F���iR�5��i�ԯ�S�B��簑�r�6�'s��C�Vyj�w�-��� -���Xs ��$��s�W�M��M̽sb>Cv'�����x<��BY��9�m��O���@/���X�y�BՑ\��ݨn�ڵ˯W�1�	�(���9��>��YYhm�\F����r���zCF���~xq��@b.k�D,Ƴ�U�[Ыw��\>>p�1̩,[W�T�)���2��u��k�R�_-/�@9U1�r>w��L����*�T�~NO�a��+_��j��T1�ۡ��w,��Hr�B2U�c�����m��a�F4~G���hnh�q�&
�.��$~�H"xd�c�~zs�@��"��#vIV�%�MC�'Z�b�V��:*�\y}8�7�����X��D���\��q�����%:Mu�U���W���ܤf+��9���ݕ��"����}��	='����I��7���c�^j7�N�Z�g	H�ߢ˭�A�-ң	Oo�1��U��~9��dLh!�r�y�W�:G4�:%�j���)7�~�����d�8�A��#��t�n0q�>�����J��N$�$��"T<��`�f_�Y͊��}�(�i�t�H4��Y�>+,�� ���,���'���G�v��%F�k"��>� <��B���q����^�o��/)�ɚ�24��B������__1	����p��}'¿��S��m�^࢞@�9��R����nv�v�G��~�h7۴
��3��؇ϻ�t���7RS�;e>��?���G�]�PH[��Wahf�M8}�:?�d~=c���b��Y���Xu�;�)��D�υ�H��~ۿ��R'��X$:;o/?�n�Tb�wH��R�,�x=�c��P�g�Y����o����+!�h��WR��)�S;؋�T�s��ܵ˜d<��ݒ��݇X�V*d/&�ZB=��A���L��E5"7����\��L^UN3.�~��y.�Uz%BM�G�LO�A���G����擉Y*�����h�nWo�`nVVZ"�k�b*i�{l�ey\M<.��C(�J��d�*�����`�:J�n�(CQd ��������E�&c�w����?��[Ip.K������f�$r�"@��R��qh;�@�������w�xҋ��u�~qM��u�d�ɫ�%ə�7����l`��w�%|��8�u�`ٚ�}��i��̊"	S4>��?Sg��[����%m;�q�M��N�.�6ƋoN)���ҋ�j� r������~���^�l���?2�2B�,���s��a�13_ ��0v�غ�M�,NU��N���I8(���rnw0�<+����м���\�̮�v)�����z�R0�a}U�����?.�i��2�3�16�9z�f{�'P�@v�P�&�������^�`@B�H�'�C���5#��S����HA��d�0�t݋�i�U�x��؉���=�Ody� ._q�<=H�¢�%�N���v �^A���
"�k��%!G��7@���.Q�����]�M�3O��s��Ǩ�MC<k\m�궹�rG��nE@��FW�(ٴ˹}���Bׅ6��n�P��x�EbQW�)��[&b��)0	��{N31A؎��h(ZS����1U�RH<��k�ͽ�O*4MX��G�j�V,!�L��O�\�fDh�ޚ���i�c?��{�C�a4P��/�m��
�Rw��j�$��b�������x��Tǘ8j�,����O^Y�Fg/7*��G��(�� W!�2�<��|���ʗm� X;���>�p���{s׷�[:ҷ(�����z��q�Β*��h�m��_�O_@^]#��GAT�?xK, ^����1s��]�~"�i�=�a���-칿�+�fR{aQK��<{P�7Ŷ$����Tǹ�<�
��	�|&��i0�Qi��L���C�<��Ikb����ZL��t-��$�����0:��^
B8�U��e٧�������Ӽ�LI8]���ޠ�g�A�f�ћ���S?�_�sY�?P ��.^!��Z�1-�w�?�����qDC�M��<'f��i��inQ�>�39T߁^�/�RkP�z�����l1�8�&��H�"� U���Z����0��7�ZOq�l��q]�t���V��e�10��O��:$�p>��In��֝g�����t`��W\���A������a��D�����zH���[{	iq.;=��^Y&����Ũ��`{V簲�9���<v��c��	��[+��#J�T���w&^�6m��U���<Fp���c�\����o���d�ǡVMJ��bW������}��]�M�¥���������k��4���~��~�8a諉,&�I�-�'��/8KO�&[�ˎ &���.v�T��� @x{�"��C:
�2|P��z���x�k0g��ϥ��?_����
���i�����d���Փ�~�R(<ʡ�����֝��3���q�gK�������u���7�x1d���n$�W�y�ؐ�ux�d9EXdD ���kƴ�B�Y[�\T�����"}��wZ����^gx�j���2fu���4��u�3�"އ��Y�x������5�/+�.8w�QC�~GL�u�I����!MP׳#�
��'	|F��eح���6I��駤���՛��nQ�Xp3�!����S�'��p��6t��R[<v����Xλ�t	qWu'ޕ�fA�Y}u`�&-
�*�<� kA�2��ӱ�`��mO���5)ЋgrD�C]a{=8D;U��7 Օ�p?�ѣn�� ��"�~�-9��c>(=gc��
hh�GY�Ҡ�ֲ��)m7��m����*�=)��m(���V�9���/����:#˪q�@����ₜ*	�n������bϾ�i�z�+����ڢ}I�Df-z+X�,E<}�*)3���>�o�5{Q��G^�~(�/<4s�m�hz8��p=�`�݀�Vb�?XG��sNʥ��*�B�����XO��a	��=����/j�&�`�� �?*nr�U��,<�j���6�k`�*_R�O���]��tƼ�Ƞ�	c��7CG;�~@Z"f��3$v����.:+n�T�Q�|�Z����3�6Ƒ������ɴ���3,mҙ3w�p��E��o�[�>r�@N��<�mxUN��>��p${��b��TNva��JNAw3�24��o�����B��J�Ap�v9���E+�X�b��B)��E��(0g7��t��ꇘ䓎N�������XR��������A�&�d�!/ ���+�����[�݄��)�s���"&+�_��kX�P�y{��f�&��Q�*���n��`oHTM�� �Cf�$��Pz� -��3#�u5R�T���F�$l���Yu�w�Ğ-ۓ�����t��107]b�}Qf�͊�C&L{�gP��5^$����I'��׊V��o"��M� ��(o��%�*���P�nf����s�/�"�p$��LDc!��68�b�^�}ˎ�&�w����ھ��+�ҁl�PP� �Q
�S����'غ̈́�˗^[���i6�KM~���ԋ(�j�
����Ѳ�`PT!�̩i"o� +5k���X9�!���C��	�R��q������W����pǌWwU��cs:T"�X�0�+d.�d���}�����PllN��9#`F�������Y!�J3� ǭ�Il����7߅�|
%W�bV� ���� ����%��c,RYŷ�3�e卂�w|xQ�K�<�}�����5S����v	u�[�I�RSELX=ٜ��a��p���C�s��o���i#��};W����=��ѳ2���M����#�)*��`���^�ɥ=�������+�n*d�0Q�^�Sԙ����$8.��Q1I��2nt�T�҅���$��s�|��4A%ƹ�I����q������]P��{P�y��\v��N�8	X!d��07�~0��n^�l��ȓ�X�F�HO��21��tӪ�������y�-�'�X��zg6�KJ�k��~+$�}M}������.�O��c�u:�Q{�n�V��V�Ԝcf�aZ*�Ө�0�kmv�bۑ����P6Ƨh|0�=�Ǝ��wң�R��Ĭ���!����������KIyB�ZYM�O�a
������'d�¦'�Y���6�,��%�G�����x��/t��/;ܯ������k�i�+�
a<�^��3�䕊�MH�k^���
ޥRv	�g����$c�[l��I�r���J�nف�٦u��O��d}i�G�xM��"�$�ϯ'�j�k[�|s�:�s���n�B�v���6�7]ysŴ�m����ٳ|�7�(?�ПfS'qR�_��;x'V~"{��p���#N� ���2�����ɿaG�9��h��4�_�ї7ܜ�,��K?A=Z��9�M��7�H&��t�g���8�'+tU�a"Tz�	:�w����[��ˤ5Cd�☭!:ۥT�a�F�o�S�P'������x�!>;�)m����g���Մ�P;S���9ca�X���_�Û�N���Ƽ����wƖ�*�M?�m����5�)E�5��e��ǚ
���3 2j���ء]v'[��L��u�e���rSD
��}�ڻ��Q�-7T ,az#2��WQ��O��k��!ӻ�� v_s�5eʎ���ng�����#h<�|���v��ظ�ks.�G5Q�v��KO�u���j@�Ϝ�F���M9e��f0?��.�b<'��B��B5ۍ�:�y��.�u?]Nd�Ll}.N_Z������\7��n� <��i@-�B�{~�M�"�çl˯�o5�a�S�����K�	����q����!�yQb�rh��g|!����vM�}C����x�O�Ϧ2�G���4�*�e���}��1�H�MP^Z��{�@��Y�R�3&������=�(a3�_�6��QEZ�B�A\6폎���:��xO�JgT$�E��g�u@�j�-��Vp��.��n�RCF��Y-�D����lk��Ԥ��Lw�%��n��n��
�A�h�ne+���n�#�I�EPjp�����~dِ]Qg���]�M��d���<��5L�]-��V�`L"�o�iD)��_�l�~�%�\��3���zhX�lisp��D�9���7i@�O��Β~f�g�/Py+���͉�>�hfwF�����]�(����8�^�1��_����1� ��R�'D�V�W|�]��SsΠ�𹚖��(�wM�6��?h�!NX0�ŶC��hF���u�n����y[����faa��n���6�4�d�;��П��S�P����Lw��>\6��g}��Q��,�t�ź�|T\&q�)	r��V�rt�ɸD�� ����@]����W��S�V������'U{U$<�7�QO�L/���Y�k9�����e���Q���)�0 v���k~�eR�ΟU�y�������9iD5�<v��G��_�'hE�<�x�Y��5���f2�D�����|�!Бo˦��yv=U���.NB��_כ9�d�t��Π2���UGD��݃i����xB��A��Ou�0�� \���W�x������zR AaR���)eK�|�Y�V8�M������Ĳ@=�8;rORs��ǂ���q��d�pȲ��!O�',t�`=&Ne�0:��U�Й��AD?Ѝ-sq+�@k JS9N-S�"Xn������o���Lʻ�)֍��D$�D��_ޫ^%\C���
�h+��v�-�r��5�������8t8���G�5G��`��m�����$��9C�"<wWlà؅ɠ��+y���P�e�����5(��\L�&���k�K�er�������.T$ӡmJ���?K�|�M�A��Dwa1L���j=�{��&��5+l~�_�6���5����u��+.�4�J+�}���S%h�#�=���h*������ ��#��#�e���hWU�j����
�{�]�W���J�]��)̈́���,� ��
��³�Љ�g�f���rބ2<T����xT�^��B�n٪s�s�|0{5���mR�+�T����r�6S),IV�L�Aa�7��2��A��'M8]��	]h�~���
۔�9��-B�����I�UZ��Z�:@��C�#Y��s�4b�Ƅ̣�H�Yo Y�󷰭A���L���Û�([�JICa3$���xNmH�2E=~P�������XCU�H�B���֪IRK`;��G��S:λ��K�MR".��J�6+���L^��׹�xLw�7���ީ�wm4x��c�Ntp�^5������K�X]r3R
����$U�n3j���A=[SC#~k@O��縌�/_�zʢO?��cCa{��4�F�Ye�"D�X�tE�K�V
[��PX<�|�cs��hسK{88�L�CG�^��(b<�u�1XG�}S�A�4��ݎ��:5����>˖c�Zl��/?�BM����uw����d����N���_-N�L$�R\C<(Y����q�7/�Ѱ�}3� ���	��6�ka_
-��-@�k�����C[��9u�v�S�SB)��i����hJJ�	-�`Ej@�J�\88�ë�W��prb�&�N�	x�@�+�;����`Jj��� %���<N���B|,�	��Q�*^���m�����	��!h����N�G^���M5�ʶI�9s����y� �xa����o#Q�����w`Q�N��Ĕ��XH\-Nǳ�z�~��B�80Ή�p�ͅllz\6*ͩ{`�}��ҰJ�Ʋ�WQ]��.g��h�j�$o�d�j���<	8�qnd���Jp���6/j.g��ʷh�Z ˥�!��'g0*�� �f��X���������<��c�.&oa^�J��p�XEkĝ��
ӹ����S��A��z�n˽���ظ-�3	��gy(�t��g�Ħ̣�٨咘��(�OD�B=Vj4ZmN%-����_��#!S��Yӵ��p[u����ߕ{�ɬ�sS��Q�5�J�!K��V��?��	����*S���L������\�p*����S����.�)b�����:������|�������@Ǥz���P�?=��ή*\�X'�1zH{�1��	�Bi���s�������7JțOd�n�"a1��[q�Ї���E�v�.SnbV(�`M��ٝ�؆Mq��Ap�kA��lH���ʈ�{�-v�����lٓ�U'G7�`����4N	�h}[�r�|X��B���1�q3G��t��;T�9G�F+�g��7;�7J~�![�[݋�F(�+뇭���9��~<W����k��J�俻����`:$��s�e7PpG!y8O�x	���y�n����&@B�ۀ�&i�4̀����'���0�U��W^�k��� ���j| R5��]D{4b�I����Icsyhwt�`m��ڦ㘩^�y���l�Գ>�y�����Gъ!�E��2U�-G�jX�o�=7ի�iD��S�G?�
����.&����3 G�/n8��X@	M ����r7Nxؓ�-2��*�~r4��Ľ�����S���V�ܕK#ey��_���Ī#&YvZ�5��͵4@	|;D��A!.L�`)�)�X�N^H;�-ҷ!(
��ޞ�yt�h��}fه�S�ܮ?���g��n>����js!�vY.�.J��:�!��*��(�h���G���ؿ��\F�2Ǆ�WSq*�7{�k5_B�"��@��+�}���PPh�����-�hn�,�^��j���*6��F��.|X;�2TIj��|G�O5�\1yLj<�WrxCXj��X�Sj]_�8W�X�e�>~��a��m���`�����C$�P�ݓ����ogogl�.O%	�N.5��"j9�t1{c�|� �� Q��.6�􃂵^��@(L;�#J�ݶ���b���M������*{~[���x}�UNL!ǫ^��{:�-ӳ���t;$�>�N�$�]*���@���Y��5'o����Ur<fh��j΄u8�����&���+����$m����H�#`.��5�Qc�$��T[yW{\�Xc�߯u`�Xہ<ߖI�q/�Xe_DY+�ã�d�{���6Hs�x`��HF:1E���b�d�e�<����%n�|)�:�E.o2k�t���*:��0b����P�{����-���Ӌ�(����=:��MfJ������@����X��i�, �;�X��O&��xQr�(,0T���-ݭ-���Ҙ���e"�N� ����4j�r'T���Y�ޠ��]VRd�3�z�vB�^AY��D�e^z`�vmE3�QK��;�X�P
|Ŵ���ς�yF�{M�� �G z�����E��`�@� ���v_�nz�y��i|C?�\<��4�.�K.0�޷��{�=����<��.�w�#*�P���_�= ��e���KKK����Z@�a�5��ef\�x����]�j�,�fG��G�{>.X~$^(+V����!y�*lUHF��Y���B9�z;�YXak��rp<��EH�
 	���^I�#�ݧ��ʄ%����#������(���?[?D���2)�O��t��\�O43o�c�U��ez$����'�H%^���Xփݶ���ڜ�A���#�t2�b'����Rt�7�C�VCA�'�3�6�[E��"���VP/d>����*HU�eK�bN�ؘ�[�Rj+ϓ��)��p
�i3`*�2w��D��l�+h�A���@B��2I�*ϠS���~`+B�f��`����UQ�]e�y��c�b,�s���DҖщ:�8(���!��!U�p�?��lHg����y�|��5L���������81AG�Z}��/��w�Yw$�li�O6)������QԺ��F���x(��9�zs�$� �Or���j�J.]n0�~|�f�tՅ#A&ZH_<�ʆ���K0�s�*�/q�g�
� ���Ck������O�8�6ga�JY҇l�6OF��R�� �4��y޿�C��0�B��3I�ESuj:@�	/`�Ù	���'r�C�Q�j}��}Q)95w�����HN
�yh��,�9.O��I)���I�E�����ȗI�i��%��é�?�P�R�l�m�������?���1*s\U��?VY,=���!��l�L�� ���/�������a���q��}���b�k�DVA�ӊa�[�$S�.�6��T�B��p�9|�1�7��Z��1��F�g�!+�n��/�.��Y��*A�0g�:�;��`�T�����|\nb "��ի�%�|_pXF�s>��>%�9SD.;�_`{�@�@�����ช��Lgwtm��-���L�7@j�c���A"��y#��j�R����_XGk1Q�κd���C�	�42�1p]���p��iӼ�odP��K1BG�z�Nm]['�������VOk�C���}���~Q蹯��F�B.�c��$�<���؟� �*􌲬�6n�]�S�^�Or���O����ɮ����qKĢy��5P^��u�j*
�;�)�k.�QY���&���b�8sfi����x�P��9-��q%,E�.@]��5�3�\3�4�?5"aAq3�8DD�fO�/W�݊��$������v�P��+ѽ�2ѽ?%�/�/���]�oc1xOIQm���ɭ��SD����&&ų�-��'�Y�ᝥA�r�{�Ird�O��n��J�]G�HN����j{1	Jܪ����DR<w�t������K(�^B���_B��󞃝����)�՘f8������o�$[�.��&v��Ks�v�c��W�&�ʛ�~���e���ke��~�D�
Y��mG����X@<�*���@+?�w���#��v���BH7��6�Xo0w0m���7��!3��q�e�Q%d�;j<A	����%L��������O[�D+�*��=r�R�,�p#Cp�z�_�2�PXI��>�5=B�h3`����ݫ��.c4W��9�.�>+�mKOl���s���F�Fr�)�N�-����R3��{��ET����T���?uF�?"��R �ےђ�}�����i���������:9��R� �A�Zբ.4�T&"����]h/_9o��;%��=�������]"9m���
WiZ%�Ð�R�|���<��V���p>�e%F�ʈ�.����_��6��w��t�t���"�	- ��w�Y��K�0_�S�՞���V���=`E䞂�nB�Z짬��?�����VwȪEDTd$ b|��	)V�@����w��N��&Qգ��%�E�� pũ=~�5<�j���g��r5%y���'u�Z�A:��[K{�x����)Q��������7���7@1�Ѥ�K
������Q�/�qÿ�#�y7�
��tFG> 
�3��d�%�����7Fάڲ�l�8+�a�"�g�:?rM�4�W����6��)�Xt1�G�Ӈ�]k����o���a�[�YS��X�L�R
�N��3��Z|3up�N�����#h�|%3)���ʒJ,%XE�J	�'��8T76J�l���j� ~k�A�ږv���y�O��Ц}�0vwO~§�v���i��4���[DdL}����v�*Uh��Cǐ�M�qn4�q��!*o���ٛ��Mn�u���	�c:s�zn���g��ل�8jB���w?zM�_��H�)�e���$�,5!���Ǻ�/r�L̕�����~*X�/E�R�b�_ת�.���G6����ޅ4^�z�� 'hF(�:����EmP�����r�9��(I,C2�c���1�ʂ2tqu�?��4tr��~�jZrDo�%A�)E6�M?4��1PG?1U����Ҝ������d��bQ5I�m�1��䤃�K�lt�Wg�g5$�P�Upq��MWR|t��CC�8f�C����ܬ��-C�	�>e�@�r�#�s���	�rXQ\�����G��\ X��@�^��<[�{���k�/bhPP��c��c2'���d��2��W�vY���(�ڲ�,�%Z�z��~��$��l�+8�ף0@�	��\C��Qj�l%��+��:�=�À�yG#vZ8��d*\
��� A� W\�,�Y9�~c�	��W�,t�?x�RKg�f"L�a��I�50m��	��&W	��C�h���{{U-褫P1}h�$��):' �~��\����{<��&5��s��O
����b	|U�|Kv�~Ȓ��F�%I�CN�|�c^�W�}9��4V�d�d���w��6�U������j�����6���'sN�j#�`�ڣ�12�r�
�*+�|!����z�)��<�8�1��ͿX9`+���\M�^�G�����9qz��o���qS��j:}�9m-Jg����tH��F�~K���48WF�����ڟ܍�� ��Lĸ�u�����A�l	�b�DZ�����Z�Uk��eV�rЖ	�	��q�zA_P̡l�����{6b.0ӊs�� Ŕ�3�!�e���1i�^���0lF[�|�7�0��� ����%,�;Tf�~ iy�DU<���F]R������l�N�
l��1O�������h��:q�-�<�����iϩ1��Ө���<�)�԰�62&Ĭk�\��ȜN1	E��O�lG��ø�y�y;R���V����K5q~�=��	����r��l&�Sv �'�f 9� ��� ���V�?^@U��q旼�e_��׿����ty~�T
�u�5�mXG�5* �T��/?�y{2"CT��u#�)��i���*X��#��L'd cVВ�vG����J��/����X/�3����y���o�H���K�)��&����!����6Zb凎ϭfP0�%���b�*�%X�n�5��2L{=y�LENW� �\�q����.m��M��ym</�gzO�!����Kd��"|��Q��,�}���U�^?߰$A���Uc�45UV�0�n�g�|��{ʹg����fzw���P�G�b%����qނ�RF+�T">�+#���4�v�B	�17����?j#�<�����-�xպH�g��$kN���V%)��z�,�+U��P`��8��̓����0��1�K�p#H��`��d|������%�e,Y�D�\��`W3x��Φ1w ���^a�$��������I4����V�\���X���7���а�)^��������
%���C-��+���N�}�S�Jl��v��7�Cj�X1���+�j��؀�%�R���gJ�ي��Z�4K�q�8����R9��#�(���8���%s��x̓P�Iɘ'S�8E�p�/Xw^P�0ޘ���.<T��?�&e#7��ʢ�zf/0o7�r�#UU+�� ��p-B�a�g)GE�te���{���.�0�j���}�Eй��Ui&�څ�]=�]=QMNȲ�le���
�J.�M0��L�2��KR��*��H7PzRi6�� ��:�8�����n���h�����Ğ���bН��ꑍ�tЂSS&�f�"d?r<���G�7���Ҡ��v��p0����G��4�om��v$�D�F�[���Z-�Ch�.�(�^�(;�/2�WC�y���C���|M��:�d�8����!}D��~]ۨ@`S��h��$�ZA��+?�u�7�p�h����J�w��P��|�X���z=7O�5@��=Ƞ��]\�T�e^[7x���-��.P/)V�rC��mK0�7���X��.0�f���"K��2���^u��?�Y��]Rb��"�[�JB]���B�ݎ�=�7g��']�Yq8U�KM.�b'�2u��3�P^ �!m��P�S
8>��9eFP�Ӻ51Zg�߉�k��{��81�62:EQ4�Kֺ Y'�y��]����.�QD�P�x(y]��*>��Khs�S��^���FRN�a�de�L9�9�U˷���fP���5$�l�O���dC�oK��w�d���Av�|�	��W k�m� �
#XS�Zj��sݤ[ªM�{H��6���uU�D�P��w(��.��^�C�E���C&x�n�^�!q(��C�&���R�o÷�s���+Hoٰ�I�e�r{Wm�v�N��a#`���n��@�-ȏ$�M�qɳ:����X��Wނ�(d�d~-�q2��>p�k� A4E3�T�F�}�������MwzX{%�<j�u�iV�c,�-��(�^hO��nx�\?���R��+���W>���ǲ�
��m(u�k�o5����yk��K��XN�$��,E�g�D��� ��5��䞏J!�����R]Eϯ^�+�{�n�C0f~6��Da٦�OY�<_���n6���Xj��ccp,Y!z?4��샐�g��O0�zb�{ȣ!�V�n���(����&����?���O���?WҬ�ʫ��G�G���,-[�e�eMv��CF��>xL�ȐF��.�K)���/�e7���D�1fx�a��:u�~z(��_�U�z�B/«�_Ύ���u��k}�?3�a�U������cP�2�V�?���gѲ��_�	���~�2h�`f+���(MÌ�'�W0��"��D��]���݋�},�556>�U�ċպ(��z�_ٝ�E'��s?��̚C�� �V��u@���b�����#9,��J}w�M� 9b�����g��z_�#M1�
��KP���!��|��Z�@Y��~e�7)��_)�_�}}Ņ���Z	"�� L�V�)"�}�dJ�"�oe��%Ssl��%�����4c�n.�F
V|��Qے�I���`����,�/�+]���F���FH��(���#�w-a��&��)���EO��[,�'��߿����V�a�'
s\.J��TtF�(y�H�K.��^xi54Ğ�6ͮ7�;%N9ɣj�bŴj̰�&ob;�{�Z#7�\��Q$A-�fs'��h�A�m�����j+�!��m�  ��� s��C�8,��Y��a���bϴ��j��Ȝ���)��l�>�*�����/��b���1S�Ljl����O�qp���Y��n(RmZ��~:y���"�������5L��l��d}�)t<]v%h���9��[�;��%�u	�n�HK�vv���o���ȵ�<�k9�+�F*���GL��(�
�3[�B�h�Ӂ�����)h�aX�FL��&K���:�(�rW6[t�d����X.|}v)��ܼ�0ypu��l������L���q-��TnAT	]`$����(Q����e~�Qc��>��${t����S��kg�_�$�9��0]�d�N�Ve���@$7�QJ��.�S������O�?�$�W�0^�:�9�Y�^¶��t4���42�U�����Q�l`�[,1�����Ik�,�����?&fӏ��yS���OTd���^�.�y�6߰��&4E�$'u���<�i��o�A��{���ؗ 1�v������aŬ_�Z�}]�骬�� �h�,��^f k���w<��M�1�����:~b�zY'�����~{ݰ�V#��<�/ � �ᠫR�Q:�B6FL��>9�Mwםd�2�H�Κ=�cd3���m��r�L�o�
pQ[�{S+���ї���.���B�RS�g��U@�6}�ܥ%W�՞��,�dk����'qdV�|7���[��h�HF��s������9�����Cـ������q�>�����'nȖ:��􄷹�ˊ��2�#^Pޕ��|y�/��7��;)�b�Q�����"ԙQɭ�K3xP;Xw�D����B`���`h�OB�Fꢀ,�M�q�N!��H�DV5<S�-M��yW�g�Z4�����~`��Ie�'c~u�\��	$����A&��Ҙ����ȧ�u��n)������!'�{`ʝdr�+y�k5�U�Ő�O��M�����ѹ��7��$���S��E)�-n��sM�N̹O�΅�%����6m���1x�۩ө!�5..�gu�|�������	y醁��3�Ԅ�|h!�i5��n���8nf/	���wZ�zٍ0
���K�w)%�9"E�d��H�`Ϟ!���-P+^�i��i��0��Yg��a��-�l�9�u�]�� K���� ��3T�b�!	~��:&�i�����ߧwla1L��"qA��Y��f^��,zaH˖�X!����O]�Xw�m�i����Z�4?�1*��'�D�60�뚉���O<�+VgI3�G�iQ&�m��}2&W.B����O�iCm�i��˚�Jt�9��^C?���f��>swX+����J�5>�g�i	�el,�I6�b�S�t��c�3���8��I+w��M{�|Tp���
�k��㭮g񤛵2���B�5���q�C�v��9��j��w�?��Y��a 9E��.P9�j@pk�Ҙp�h���^3�	��>c���S��͛�D &vIC7��:��%�T���VI�Z�V��"B������~�+*׾�膰�@����ZT�PB����5`��X\dR�p���QР��7�:N�����n�Ԏ
�PQr�@[:+AuiG��� &8̾����Y��r\%��=�,ˊ�>��ؐC
z�S�Dڛ����r�wY�F�n^?��ߟ�c�Xs�]��k��Adʼ��`��D9��h�@���M��*L(t.%8�P;|��֡�u/���"R��+�dU�.�`X�=<�$����Jŉ����6<8ٰ��b��>�5�lB����8*�א9�`#���,����RxU��9��L���Y�V�q	���y=��/��|��J�Lrd��*����� ����[�Ѿޥ�H�5Gǰ:a���<՞�Cm�s(b��~b�0C��Fk�ZdF--����5c��n�`rHV��F;ej`x�o�}�*D�iN��c���Jk@���$t��L�qZ�&/�B22%m:�O	l���;ܧ�J�6O�^1n?������ܼ���ơK�	t�z�#��Ǖ�����_$�r��y�A(�z���$Jnw�.���v��%*Wr�,�B�Vy+���~��`$X��@���o��hv��+0�6� ���4�rC��;[�[���U��VC�p���ɕ����z31�O�J�)@L�0��v>��n ���I5�]� ���N�hT��V�4���)o6u����%5=�KƢ����l�酂�7�B ��xu��K2��_���; �uln1��o�|�5��A'�ދ��K%�xxs��[۰IxnZ�s#&������2t�X�?r9);�)�|p�R���N����;�|���C�͊� B���Bt�ǮI�X�8���|��D!���i�Y�\��w��"B�sŴ�87+����3P�j26�!�Q�c#k��� W����c�:N�p���ś,�?� ���-&�N�`|HE�&,B�L���p�{�^�<O���e�������۫?VV	���IG;�_�m+��j?�4X"_&Ǖ��I�5-�ϛ0���!���Lv�J�цA�0iS��f�?A�Q��'y�����IO���`�|�#lل&��:��t놓Z��v��G��뵢��F�|�T'DL��5d�Q�}�P	!���p�C}5Të' l��Ts@��(�	���-2���{is���v�ߩ8�ѯ�TvC'�:)6���+6bfd�k����zS�R��=�P���u��X@��1�5�U������K�'�c9V��^���Z���9JQ1@�֔-i���a�"(:5#2�*\�&<O�X>8_�z@��*�W�(��a�w�W
���[F>��N��g�v-��X�^��}�E��h�������{�L��H�;�!�&6Ն;�:<����FQ+7G�L�BkeG�qz2�cΗ
�G���9��G+6�	��Tˁ"��U��)MTz^���}1\9;��"/�����l�O���<��"�Sj��w��gc6���[T'�����m�����d�	H[87��#�\����Ɩr��'x�a�6�Kaj����jE�����u�M���n>ճ��N�7�f�jW�O�K�} 5�B�%��\���G�m��]�HX����y�5��)�@�Leh�P��aD�%2�(�
x����B�A�<�t�l�O��z�y���d�k�[��A#��s�@�K����p�
٘�.SQ�[��gtPa����jn�W�@%��: �Q��'�i�d�����l ��DB{Q���e+O���#khg%$�o���M�.�=x}���h�sP��5�\EE���v�Ąw�K*E�ɱ�W�C�T2���x�Q�{�bK�<	��r	V����O� }M�Y�q�9��"���N�+M�:�ߣ ���44�Ax{VcI�ݱ���Z�Z؁�ܨw�>$p�[��RܧW+">����M���C���A���G��X�7M�F����*��Ș`����O�ݦiZ����y�ϭ#��P|Of]#rӡK�4��OT��qL�Yx���)dNR;�@���
�L#�K�Y�N)��D��8���BB�s�hc�z�KU\VS��wPؘ�cU�/�ƙ�49�k`Qn~���ٞ�h�} N-ǟ�
���NIRw���H�Y��yhcW�篤����9��j:��c�Ї�k�^�h��@XE�%b��6Z�lb�=Y>X_�fKS�[�hh)P��~#@�Z�$oWu�xM�����y��fa%������}sJ�hb�h+��eؤ���N6��8]����U�;����r��9�(�L�.Z�$Z$�o�]��8���Ѡed���0�J�+:n)ئzI|��&O�~�j��\�4��|�x�Z��U�����v�N�(k�-��Jm�{9F�m d�Gk�G�۰��je�`-j����f�bˆ�@�}��+�VpT�f)��0������h�d��	���0Yž�L�-��z�u��n�B��O���{�O��}��+�t�l���z����a�V@����5�gl�喭^l�}�o�*Di�|�cۥv��a|:�_&�$D�t�(7��|�LwQh#ƖC�*�R˸zd�EQ%1.�ƹ�s�}7J�4�⑻��ڥ��&R
��w����M�_6�#��޴x���&����~��q��ol�������1ֲY��	�U{)�o����~����W���q�D�5z>�X�,������G[m�,��̏����UICD?�����5�D������������ڸ�X<����_0�g�JH�-QP�SM?�$6"�a(۹Y�|�C�Z�4f?!P�-�b� !��T�%4����#s���� �[jh�h�*����5w��$1G\����>c��NQ��=A�9<�<�?�-�Bdk�0;�W��)��EZ�xp�IC~����K[�9<�	-�}$&��?�k����"�ph>�IV��6� ����ܵ.�]�A#f��p�*l��| �#ڶƓ��!��)�V�9P����D,�খ��A�4�� ����.O&S�t㍰q3���=.�ha�=O1�������2����n��{��i*2��{�:H��"=:�2�z�gb�mĿ�3�����7�G�ސ�s�G�*��$d�.��WG�n>g�Y�oY��s�@��+Th<���2JU�*�ʬ��v�s�Y��j������b·Ov#	j�of-]�ȩ�w�mc��=CtT��NS-�H"��Kȹ����@��L*��3��3"b�ayǨo��m�/m��ŧ��|��r#��wދF��ې+8}Kn��يLW���Jz�Y��u��Vg��&ypXU�nkt4�ҡ&��*���"ԡ
��Q9�"�L�T�CR�`i:?$_*%9��w�9�حx�^Y���XnP@�A�j�����_�����!S\��Z�H�$�g0�h�VԴ����G#��]��[�����(�'UbG}��.��:��(�p�IZx�"���	:���YBWRP ��X��P|� �d��|^UnU�8i	���d��o�;j�6��	�9|�����;����aP��\����s�s��o��du�2U��?�o����茛�s8u�Ó�X�^3����b:�
Ɲ���}��Gt!&�	��(� ��硾��fb�i[�����\Q4iB��)�n�:�F������F}zwf1�]~��/�R+lE5�� >~W�TA����ntE�ֹ��Z߼��m��7
������mM�+/�wc��kP妫���Q(����;�z$�I�+�\]1^�R)�q#�����s��/~�S��
S���ޖ̸~��`�Tq�+x��-)�t�20Q󵾏���5��DGP`$��a�6}�1���d�Cڿ���z�P�&���^#,?v9�v�(��ny�&�~�R��19 ��� �X3^��.v��D�|zlg�ԧh*��c�$�bE�o�|ղ�Bxl_NW��rg_3� T���0����ܑ.�"b��W5Q�o��ɳ��oY;c3������I
.*Bnf���x�&��鱈L(0�K��p~,�jص!�ܼ[��qC�=��Cq
0�~S�~�&�Xy�C���\���d�����ey^o�|��x��Ln]�3�F ��7ǅ�ϐ�x��=�������֝�x��>�X8�qx�[�Ov¼��'��C�-M����ա�����Spt��.�ȡ��`p�-�{��i#��@e��*�o�X�n�t1pX�ۈ��i�,թ��efBlG�{Uڭ��2wR��1�ׇ�̏�]�8a�<�+��/��W��[+AW�ȹ��s�7 >M݊��>p��ΫL����yǗ"��c��[�w���]��"�O�t��'R���;Mw�c:4:���5䋷�
.B�z��B��(g����ǂ�XN'3�4``���ФfǪ�@���7p���;P�,�d_�F"�֎�4�m^�I+������-%*�n5�C���&5� �<�r�3=���R`(k*����g@y'�ΐ��+iqju`yr$F/B����R����f&�}K�ʕ�OE��-��:��� �A�}�qV ��މRgH!'g��F�Q���^�<��3r5/�%k����r��e�a�l�.\��d��
����Ҹ��8��f��h0�P�"`���7���L�_�.d�
�:�-�+�jܚO5�M������~�=�]f.�����W�-(��>�G�-���`������^�;�y�sݔ6_�Z����%,lX�#{� 	���Ǚ��j=߈��J�J~Ii�s�'��w�p+;���z������C�߯b�1�3�Y��� D%Qz,te�z�a:�%b�"�\b����Ff{�)�do��A�?_;��n(f���{�aJx��y��᳦��l!�9��䣰���䈛S��_LNz�z��(tl9�V��>wK�����D3�ॱ�l_�'7�ՍN��Ogy8�R�� �Ԧ�NoR%��k9���׸{&ѕE2t��c�,I�qm���Bm�.Dz�d��U��ͺ�
K.�և�B34��H4�p,*CiW� �Ǎ�`�����/��C�?6K���'O}d		 1��t-��_��՟\�%��q��t^^�T\��0JaMM�������86����x)=5t��*��O��U�5�	��"����y�ep��n�=|px���#T�i4"�%h��;���#�W�/ڬ.b�E�MX�M!2�q����j���p$.�sau�6 &�7�j���g�d3d޺:��b�-����E��8���Y&��8�I����%�����.S�y��ϊ��@��Tt̃�?�˫�� AK�bXa���A�p3��p�����5(�d��f�`���C$�Ҍ�ȋw��v9�T^��pGU�po����n���A;D���Y�C<)�u�znwԊ�zK�cK� $[~H"��}���u�����+�!�q}f�"�2ڜ{��*��N���-2�Y��	/htd9�K�vG�s=G_tyEzm��8� :\<��RN~XW�_ǀdSX�j洍a!�o�O=d;�ߜ�t�wk`��0�IE8��<?���0�ߚ��I�?�#2IY�"Zqd���g����U^���BL���9�%���AS��$��Qg.:��w���I�^���A6%�T=��tɅx'��N<���u\�L3�)m#�Wٻ��s.�|D�XТ�\�D�yǱ.�G|c5ƭ��/���&�Y'�.>�T[����q�qg��1I�d�aX��H~�Gጶj\ִQJO�8|4<�*�"���`��@�����<i�K����JG�9 ��q��N���T������-;񈴉t{[�9V�<n�����o�T�;����i ���o���$҈T�O��r%��_ZD������A�ZR���cx	�΀RU�\�GR_rJ�`�ө~��S�G�)��R,��[���ȎqJ���Z�ԫ ��j�k���~����xSs�-��=��$Ly�����K���v����U�㤈]�&c�rA6@��VI�
j9"�J{���c���i���l��R~V)fF�����^3��ű���-�[@���ƅL3�q�e��Q��i(�Z�_�	$�o(Wu�j�^T)[�#���]����h�4ˑ8:���J6y���k��q̅p���X0>T��/CX��bE�#vVP��Ĳ,�ʿh=XEƃr
w(+�%-�J͙m�����f�Z�iD���h��N�Zo���j���
���ס.i��z���ɂ�al�/0��޼
j٪C��V�m$��kk�y�K��lO5"_Y�A�|?t$�o
��y���bYB�����-I��Y�E7�E�̾��O�S�$k�M�m�]gq���/�Q�ɇp D��nFKe�6ʧ@Z���k�������I�.�4W`��b!Ht��Ǐ��w�G�!_fQ���SN�zp���\�|t�̉���d	2�#�t$����7�;P۞:ØҎNl<@i���fы����i�����?���?v2析��LT�֨K��4$��ތI�⬜#���V�?�Q&�B�K7���v�Cj<M9�"���,�
i��VKP#%a����Cφ��a�q�?^{����x�KTL��[���tԬS��o+«`�pA��N�zAy?�Z���k�������U��H��+��uBߺ�,~�t&u�D��1Eme�U�U�(=���!no��DC���{6���n
*��f1�ݺhR�Ľ�ޒ�o]mȲ��e��Ȯ0����U��ޙ���Y-K��Tt��%��&����Oj�����Ί�U��FG��/�Ԛ+���XܷV���zo'��n�T�#㐼 �ʪ�,ebj��<3���N�-��o�\WC�m�Y���RQ׀��:�,�G����,�e$������r��kA�!Qؤ Z����[2;��~�K~8肟��u�T�X�>�� ���=��~O E�������.0�o*�"��v��ܜ~T���޷�Ű�/��^�:-8��o�♗F�-�;2�1Xgq�*�9�^Wb"�\��%�zm�R@74�y�%. �W˜J0��G4"o�	V�N=��K+�zi$[��P�l�] m�P��0��p�v���r�3&�S�׆g�o���d���̛낦.���U$�hT��k �1�U�0��e�ܙ
]�d�N5]ҥ�Xj�f@bdz�L(G�d�[[Fn���"�1.#��9X�k�.5�i@�qO�J�u��9Ey\�xV���%��d�D�ݓ�ߕ��5O��1�T4� �xfv�2���s[�q_��!�I�,<)ƛA?/0�7��<E�p��­&�f{+n�����L�o�$(��ȧNV��N����?D%׶%�N.���B]��e\`x�ȃϼr��3��$�?�F��܆델i.@=K�.�Az����ߚ٭	����� ��j�:�X�2J�N7pAA3�ӞQ��O�����\�$�,�W� H�$�L�CGGy
�`r9 Y��PI���q��z��p�X+������#�'$H���2�0��v�>[I� F�z/,��tuf�n'�s����u���o���@S��ɾM�\>������L�&^Ve�n��P�R��d��]�R�`-}�b�`���P�I���ޯ��(=c��I����ӰC�Є����sM�xi\E��OS��*kD�>�X��IS������0���ք9P3�U�߫�BD.�ֹ1WL9����f
ݵ�:d�3]��?�n����PЭ��z�Uw�Z��( 3Y�d��˟+'�f�����	��d��D�s"���u�E��mݛH��Z}��u`�a"�|Ht{�n���R�g p�_+=A@>�2,�Q�B��l��6��0n*�Vܓև��S��E��!���j�y��?�4 �3��27vK�y\FG:�~@8>jH��g�W����a�UoT�c�.|�+�!M��f�s�䔒�qm~��H8[�����By6����dǅ��u��[&mf�l�k�]ԧ����M̔��e	�4k*Ť���ɾ��C� Gc��L� !�ٹ���/�x43�w��HCc��%�b��"Ϛ5g�j�1�pū|��a cG�
�7j�E%Q��۝�y�H��e�R$����㝮��W�_�DÁ��4����H�or���h�Ѭ^v��CWnNjC0\��ʜ si�FƔ��q���QC�9Z����W��U�g���a�Br)�t�ce߬�)�`O�aAC7t�h�&C���}Ѻ��S2U D����j�'���hNs7�%+���T�D\�������[�$A�nV�%�d��[^�Љe���$h��Z�αj2����%�x��m�K�IiB��-> ���Mu���k��"/""8�	oS��6i�U�e���� �~����F�X����5�� �&B��ԗa��I7�IJDj"���TIA܆���?����T'������S�V>����cO�6�������m��t��p��C��p~U��
����'�v }�DEv�!��Q��tKa�)o[}
E���!H����J�n� ?�dqp�9�D�`~DR[_�YvV�b�_�絬�"7��6k���R�\��7��P���Gbꗓ
 �r����ǣa�XV�
|m�����@��wԖ�r��&�B�X��PX��Ӥ��7u|��J�Q�L�"�#\����Gew����`x3�m;�$�����373��̛�2$�QzNr�Ғ��a|���	���`�M��n
�����;cl��6{��;��� �lr�`�A}U��/u�8<]��/�J�I%)B�'c��7��3��I�9�����V^�X��jS$�9��ى���ȩ�/g�o��:�/?�ۭ�K30'5Mҩ�ޡ)^�]��F��XO�r����;_�.�>>��nlIV����𦅜�p��p�+l�IA�[�ݙ7�����]3�z?�=O�c-��ƥ�Z-�׼�Ի ��q0W�A���}2��q���@KҲP��)�U!����2D�B��s��Y&^Yg*\�y�	ቼا�L��*�6��ʷcn���{���ُv. Ez	��c�����r�
���DW6,_ו$�o1���/{u��9��]Y~p.\ʽ������i˹�}�j����N6)Sl;��1��X��݈A�Y�O�4��e',�j�y'�j�y//M G�]��N��L  YJ{1)���M���h��L�t� �Eu���$���՞�&����,�����d~up����:
?�(���}c	�;4�d�#A������.z�e���~��ݒ�/pt�O�~�URP��}�$�|�$�߅�]?��Te�2�VEoSh�#�|�!y-Is�c����b��n�S���M���R8��9)������̞�QT��Ck?�p�� ���D����\���h��GW������`�8V�w`��w�7�i	=~��ʲ��9E���aDJ��1�%��DM!9���n�����B�K�.��M��N�Ƿ���P���5�������.�϶�p:��1Б7w��^3yjec���n.��5vSD쑞�3|��('����#-8��~W�����}�����֞�;_��O�[���r%X��{�:��s���<��l�?�7�P�vC�Pj�!&�U����e�~X�1�,R�u��x��
H��`��CTR����eخ徝4&8ѱӟ�H�8g�8�T]�3U� �A���^ֹ�44�r�.�r,S{�8���6bR��+{Bf|z����$Vd�N=�b�pm�.�=0p��2�zxO8���.�
����}�����	�Wиx�l7樉PM۔��'��l�[��C�Y�*�ݒ@.�TN�$�ߺ�:�.����~H6�J�Z����~Q�6��M���{2��+���7������0�M��
 q�_�-JwW̽P�]�R���Ȁ	��=;F�
}�[7LJ�w<)9}`�����01����Oe��yb�D�j�\Yz 1�j�ܸ
���8��� 멜4*�-�������U�X\sO (����?Z�)a��I����R^Ҋ)Fw��e�T%��z���Jh�J9u�R�K���或��]���tʯH#Q�h8YJZr_(���������Р��|�}�4tj &���n!�@�j����G=�d�}���!�8�#�q��U�*�����`C--��;�{��-�)����izŨ������5&�����<7p��;�#�w��L��f�M,&�l6@&�s������!T�c�t��Ů����KX�4q߹Z��� ��>Wh�t�*�}l��m	����>8��� v����@����@K D�7�Gn��`���9W/k�j��>��6QFo��u�ƍ��i�U����"� ���fq�~��ן��w:^(��,��;�&
qLڃ����	���l�Fq���i���'���ݢ�$��l���	���7(A(h�sؗ���%���7��t��0�I65]"��	y%g�ǘ�ev\z�>�iU3�����",��GT���<=`�Sc�]c�`���x�L�ל�b 
t""��;�]���UXU�
O�"x$�qS�Y�'��)>��\K��أvn�;WC&�1���,e�͞3�Qv�aO�Ś�^��q/�]�ҋ K�lX���i�(�ۻ?X'�ߛ�S���A��1_ax�MW$�*���X�g�#�
Z�`|`l�cŚ�Ywk�|�\_��a��T��z�J����L���9����İ���U�����/��>e_�ԩǂ�0i��>�y��
�(>�
DY�3����m�-��SdW�-U��%6e���EE���X(�/��J�3>w��"\�W9�F!f9Ͷ�q�c�G�'��c̹��ۓ%�>���7���:K!��*�Y7�*�%qe��zԧ���~���X���"�gk�����K�1����j��j.�I����!ZU?>�x��@�j]=�~Զhckc:��@D��5��{���"�S=G_W�I�U�yz+���O_���n��a��$��Fc@S����g��?E�a�)�^Tu���#�\��q��J�a�r]������x���K�����x��ߍ#Y�-�zY�	�o��Ff����WZ-})]rI���l����2&w��4|k� 7æ�}9 ��&,k�`@�Xj�C|{_��,����d[0�(~�[
<`0��ڨQ���#F�+��-68v,����M9�mTj�7�w��8�7����7!4gy4�9�uV~a..���R�w&��.uVi�ħr ��c���6#gȁh����1�K��m�K:��J|�וּ��N�HD�kdi�p�
�_̙��^۳�2�
1il�X_Z5��i�m��L����\��� ��w��B��V����\y0�-e��3�0�}q�CGC^����'0t�
$��V<¶	FR�;�/ņ_n��6��NR�p+�LΚD�9Z�m�W�^����pE��#7��,��"3p'a�����(���
��<ڭ_p99����O������K3�مV���K;/h����Og�z!�3'\`��$�"פ�,w�J����v� ~�DV���tB�|����`peW�w��ި���pTΛ��#>���٘�EgU�[�n[,K��;g�?-��z�on��6<���A�61q�>�rÐ����
������֞i�3��vQ	I���	h��-��S�0wU��O��"�� .^�`�]KO�S�)0+۲R��,W��ޱ�]���¡(1���QT+z��4]$�h�Pd�M�����[��e��Qd5ɡ4�����.�*O\�'REݳ�ۼ̻t,Y�H_H�y���6W�S$v&��������:\hW��U�5U��"�g��E;�w�� �?�;��ೌ���-4�:��ޠ��9�眧ϊ3+ӲF�v#�tx~����UO^,��;<ry��*b�[�#���݃9�Z�4�Fh�[X�H~U#%(��� �Wv���D�oV���TS$��r�uR�\Np��	��q��h�KS)L����U�+�w�_���?��s8�3>Q-^����uq�[+^qz�嬺�������â�2±��.᭽Z�`��=��{̎������NĜΈ4Q��ϳ���<����rmL�w��!DT���-'3Y�|�1�C��O��B�L%m�4���Up2`,�Es�%�ͬ��v��u۷M��;�0?jd�ܖ'�h3$���']��DĠ>;e@����<Ź��/�
'N<%k��P�Kz��Z�,�f�f��@�$W�*�j��J�ߤz���/�!�e}��v~��ؠ%,g�L4B9�e��^@�oH��I�Z[C$��K������6��;�Y�iy�KF?�`�냒im[�2$�I(����!��]|�@��C<��XIYW�����$�y��/n��m#]��w'%N�v9�"UJΉ�~�X{~]��dS!��4#M焇�c�e�ż��{�u�,Db5�4�_�+���y#�^KXp����;m��$UX��N&W]�3?���[���b4�Lx*U�=�*�Bg�W�	V2�ȉ�1Ǒ���p{��g�f!�	�|N��B���2���^�J���|w�RKlae9�D�.L+4�L���B��"<��	�<�J��'��˨�x�1��#WI!�@!�@p�o�e}��K�ʩ�}w>�U�}��ґg�"�&<�2)��)�B]�Čy�׎�1wYGͺ[��r�`�K��s�\'2������%[Q�d����Ņoks�i(��#/A�-;�H�~���m<MB`�!��~���8�d؄n?�h��I�]�ZN�Ij=��8Z�-�����n��P)}�9��cE�� ��Dyw�㉸�j��<W����ц"�I9�����-ϩ�.��7%\K���roӮ�Ikoۈ��Vټ6�a���#�LV��#�9��MK(��p��HkE���Xu��,�j���}�E`Ah��<1%�ڨi|hL=uLў~�N�6kS�SFS��k�`?䙷]-�1r)w̂AO�'�G*���B��1ǖ�5���Z�ݑ�v_�n�mm�LY�6��㒜�=�'3��?��D�]���p -�:�9G�a�u��n�LGS�^� ������^�[��/[5�4��"=T�vp�!
�����j�˧h����X���K�"	w�9u��5�e'6'���c�꭮��{'/�`�2�|�� �~w��gA�Z�Ds�*5�t����ꅫ�{�KM��i]�ԁt,�r�!T�g���8T!	K_ V@��v�y�8��A���6��*���zK���M_捛�̪5~?{���$"���og�J���	o��̻	�E|��R�>�?��n�\5�׆ڪc�O� ��U�O)��;�+�T��0��s�b�g�M�N���a���&	�on�)���H��D	>�'P��~�ّ?����F��U�'�+>/.;�I�v�}]�tJa�3ƀ-w%{h!e���}�JD2������/Jd�by���'&d�F��p��A���<E �ۑ�����q��Ư���2�Oҍ�È��:����-w�A�n��ș)�T_O���/�p������4�G�����qIQUGA��8∙�n����j��d3~x��:U!� (X�p��I�u��6鮔C"?\؈�[�޶1�*s���0�e�{2�����9X��
�S��|��k0P˘����п��^c�" ]`���G>th$��0LY۹��SE�a�>�ʥ'�ȏ�{c^u4���˶%��ԥ!S�Mc�|S�}3%�B��\�Qў=|\Rq�-����uY?DSw ��Q�e`��_"+Ǟ�DN��t�S�Z�}��a����P9�y���ǽ��CMp{m]��z'�L��&���$�05t���t��b�w:	�H9��Y+�-��+l#��	SD�Q�dNF`����~�в�?��u�fHq0�yn
���:�8��/x+;%g��B�E$���[�*WQ�=���JŴ|6������bn�{�-����W��G�E9|d�ނ�'�0�B�Ŝ@#�֔���>Q�Cii�@���n�X,@?�g-Ԉ��{u����ާ�W�v%��:"�ɦ��Lc������+�����e}� �}Z�q�Ĺ����ke�k3�lSJ��u��A�Cuԩ��xr��3/&Ǳ_�������F��)�d��߿�H��ft�;T̈́ �?�YD���w��͈���˝���&��N�V��k���?�{H�m�O	����Z^�cE�/?������~drg_R�e*�d@�C��Ÿ��6 [�4E�]A��٘d{��cDc��M�pmP.8��[Ir���55Tfl��J��c*��.�'9�����qd��kY��_��Z ��Nl��I�%����Ǜ���N2�	�7ȹ�a�Y^a��Mg ug��0;s.���5����cr~��D{�r�p9���4ҙ��5�iO�� )���Kr�~c�a���c�^��0����mZ���5�����B>an�ZQ�ǹ�D�I��>�]X= Ё`ⴱ�a��}{����~2�#bC]�PC��v-f�w���-�趬��,�����7�.���l����6�1�s���_��k�e����M���r�8��]7�e#�J���s�-�Yk�|hC�9��ԣ��+��Xu�k����~٣5�6#C����Jb��J1�9x����Q��������rB��w���e8��NǕ�=�55,*��h�7����u
�'�qU[�%��h�2��S�E¯�;�@�+�TW��RV�v��g^LI]+#�d��Xa�~��� @x"�>��N����ڔ��S���H=�A�n��ĕ]�C%QrT-Wua��>���k�ʫ6�>S��\�q�9��R�σ�|/�B�ڪ �ԛ#�l�U[�����Ŕ�A7�����d�j@��b]^y�2�Ŕ�Ⱦ�Q�7FK��E"��ǻp��&��]�P��E (aʐ#��[ªL��s�k�� �)8�!<�����G�G���g}��5Up�쫦�(���5`Z�s!�5Oϳ���Ʉ�5N�uw�q�.�0���<z�_ݐ�X��{����#�dQ(����Xhr7�E�^�gb2UBNᚴ,(�HD�J�y[;�{qJ�?G@���ӵ�*�u�R��=��0�+Y<��AO8�ِΖ��?��7K%	,t���^�Q?��]�$���% $����5�����D�Y���$�=;KZ����S���Z�D)��Z���|���I����G�,׼�2�:�D ���ħr���.�JN�B���&#���y�T��5���N�tA��rr��;Q��Z'c~�-��b[F2p�*��<�ݱF\:~]y��|{F@Ld@d6��FlOs��dOB�]��BĦ�j�V/� }����+-S��XJh��X���Z�Kܰӌ�S�\��ZZ�sPh�UKH����ɍqc|�h����3�T�:�W������M���A��#n�R)�X]�7�ly�� ��,		�:�%�8��?��L'�C�H8�i �r����Ŝ��0��+\�y�^����%���N�4EFn�C⅗��5��('\��a�����u�i��
z���Ǟѱs�rvZ�*q���~����_J{�ZL mY`D!�bg��N����m�h�.2ڲ�4ùj��!]"N���؜3�������>,a�_�G��䏜���h��Ƚ=+�,U?��A���&Ű�d�x�?���X����(����-*B���������,�+'ө޷�eV�Wt������1>@e��Up��t��$9aʝn-S���d�-{\,�����t0G.�cA+hz:ƢV�i$�"������[[�M�='4�}|w�p����/�  ���Zs�X�{z�ڠ�C���q��@{�\��y�6֦��OYMǐ�b�*�'1� ���v�ύ�o&�PN�j���a=���?�^�ʾ�6�3��L�dn�`|�͗[��yCέ̼��?DzO�jjC�p�q�y��[�M{2s��%��LuDˉ}���W�Dg��rie������s+�{"%W�Uajņ����F��`�P&L�gd?�Q��c���1�֯`�����S٣��C�م����4��C9D����d�wr[W���J*�Ö���j�n�cN{eXX����7]���-64R�Ɵ\P����_�G|ɖ:_Ϣ"J��vZ8�â��2o��C������5P�/�CS��;��.�L^`h��&ˎ�$*HvR>����%SK�q-��g3&V⫶vZw�T�pOR%�<���臏L���̣��!�x[9�7Uu�v[°1 J�R{8��F��#�Z^pzk>��f:2��ڥ�b9Yzn���xu?��d#<C�=�m@���~nTI���:��sl sTb�A�4qų"���529ſz�]&�Z_z����'�rl^��v�a"3��\��5��'Aú<Θ%��P�K�i��<|����u�|>�������"a�I��(��<���j���_u��Q�ua7(_!��i��4z'tp���')>���`J�*��<� ��&�RwK;���ӡ>�CW&|�>�����O����/x�M<�����>����Kk�v����ٽ��m�G��o9y=��[溈�����EYt]c�*����Me��j��$;i���U�H�s�R���rb�M��g�)O�A����8x�a݉CK��>R(�?a��(!��pC!�)�]�DIq��^�����6�i�017��^��"
�	��^shQ� � u4��X��i���ŵ��2?c���o�2#U�6<�!�AjiYr��-�q�$(:�܌TIbg;b*�g[;�t;�s�s�:�x1>���K�X/�u�?�r�g���O�H.!���p��Y!��
�,����\ܼqiP,�>�~.<�'�C`�q�
Oy��ec�w�Q�sB�A�Zh'��)��H=�M40 �$�s�UF��W�a� d?2�~�V6���ťk�në��V%��y�r>]�T�f)���%�M���J��o(�i{��n4Hn�  �4�}��P�%�C�ŵ�˂b�*J	Ώ:z��5$K?��)X (=	q�smA��Sg04,.`~��tJh(���_���pHŘ���ۃ�O.�|YW����ԌnЇd��X����s*�t�r�+��H�^�����SG�`�v}�	7�1(=x<N���%�Ki0I�t�'K��|�a��G��هh���D�G[�ȈI�~\��!aM�����2���:��K�����O����p��>x@Or%�s��`o5�h,t^�' �#���p�z)0�dPi�����������!ZQ�}rF�}2�%�a��f�Ch=�T���a���� �[�o��K'����EK:LeQ����Qw�h�ł�+�PW��ɠ��2��p���7����+�7]��%M~y����!x5g�o]�
GA�]��{e)� x�aSȈ%#`��a:���ݟ� ��~�Vhh����hg�/��$˓8��s���8'�W���.�����!����:0/�Kl��1�;s����ib�n>,��A���jV��̸�9�t��)~A=�x�L�Ҙ|yy�{�=i���	�'����E@�����<�_�±�G;&4@��Q|;A�Z��d#g��+������ڟm5U��Kп{Qm�NZ�^��o�~�U��X�n}m�	ж+z�e=�u:_�]�K�+U;��>�|y�K����KRN�1��0puؓ��W��S,�Б���:=��D�Y�|g����G��ӊ�ˡ��0�}�S��E`��̈fy7�"���j�"����5�������OuEH����,Y���K��S�� �Q�L�tZ%�/l4���g�	�#0§?����d�Ҁ�J�v�1T������1x�ܜĔ���}c����5�K�����P$�A}�xr�Y��	���>۫,�j��z��� sn�.5�&dH�~ϒ�T7��9-ĢA�M�G����O{<8!C���Sܪ*�����<�L�<�8.O�>z�^�����T��r8�4�W�^�@$UK���M�r(���?�s������KS�T�xAI�vS��	��ypKe��΢�� ���/AI�+ߦ�h|��W>�����E؅�L�/JV�hA4���x}��r��l����mk�7��>��̊���zE�)-�h�P��B�E­��ނ����[*Z��[�%���+��2�}-�઻*���0t����ēb(��n��f���^�G��<VK���z_�G҅a�\SШG�h���RO�ز�f�AC`���D[޲d�a���l��*�MS��P�8��xR,�F����!,A�0�Ca.'D����n'';��֏(ݠDE�C�.W h1h8��ۉ����N;���&&y��Su��4����g �WR2�U�9T���q���;�F��3IO"��ZK}�@���T�c��emu�nc��F����	D]�[9C�;cIz����|�W���g�:ǣ=�'�1Y'�5j��D�������oT�����<7F�o�>(���ͮ3BY�a��#����^�R)�
52��"�g�Z���p�O=�Id��yb�����X�o���Ka;���y~��:N�T ��,�7Eq�aNzv���1^<�����X���8���7@W�j'����ҼX��q�Y�f{lG3a�a�S\NN�\���t_��!�~(n1!����jo�F9�m�p���2�b�[�
��A�OrCY��A��eV���a=C�.o�S S̬�f`.��_�r���I��}ǟ*:��ꆱ��^�+�1l����3����;+���c��!W����46��4Ѕ.�g��U�#�3	2�Ia�JE�L�������q���E�PJM�v�	0\�+�n\���{U,�6N@��F��9��7���еtK�0��RA�f�#�?^��ê (�U���x��Ư���~��wޖ�}�'��K4���\I����?J�H	M,� �0�!�%�F�a�!�e���e�U{��]-��F�;'�փ�����KV����"��=&�x7s 	FV�ߩ����5]����ጒP��	6���/s���ǯ&9�V�Y/8DrfG�Ü0c���U�ngм�P�{��z��?ӓ"��D�_��O�6}��
�HQ/���Cp=m�jG%�u̧씵�3uB��2�L�X�i���m,]�n��+w��=v�/�&�"
0�����A��	�Wkv�r�
�j�5��C�ߣ�o;��G/	�l�2���>��lMC+g����4���:�gګ��m�F)R�!ß%�g]�E)G��&9��0��{ ��k�s��KYG���(�K6a�\������b�7`{CsE�����t2�����ݦ::C(���ϰ���%���+t�3�E�l26��Y,��FN��gvf��lbl>�w�+�VW���!��>f�U(L����J�Y1�@_ޏҦ����ՔIY"	��8����>�pA5a�]��sj��b�0�dx��+F�w@��^l,�]��x�e�oj��Xn�O4蜆s޿�S�ϧ �X�4�=J��3���u���-�������&�H�1���]F��9�-��f���Wa:��>�8[W����"�e���tfLNR��S��=�dU�ꜚ���}G���w{K�Ml��E曓�݂)������Z��ϋ�`�Ή�9��,Mo 2a %�)d(b�0��ӊ#,K4C���@<�oNz�����\�����?���&��R�"`��f�vZ߹?
_���^a���lND�8�*�MҶ���&ǔ�c��/=z]�p���&o��K)%|���#��QFX��l�!'����S������R.nd�KՃ��d]] 7���Uk�ƠD�r�����:⛱-<�!w�?b��|>`0bE�Y�W�׋h����weap��� }a)R���1���u3�V�$g�8}�#]����%8O����Xl���,S��{���2��b�]ha�ؗ���O�����A��Hn���M���Xd��#1Gf�Ў��3V\0��)c���\��Y�ַr�#_`���)&}�OJyrY���@)�
R
������y�˿f�&����I
C���e��NH={������Rx����)����)���h�d� 9"V�����c��W�P��5�"���.�6��PC���Z~L�3U��0�R;q㚌�c�ص��T�>A�𬬥�a�](P�.�4#M�)Q��Y�<hhw�ت���X�ya�]�H�a��x]uE�~����1��Ӓ(9}�<9���n
��Α�� ߆�*j���p�������(��I2��)D�wC�
P���LS�=Ȱ%�E����./�k�#w�܌#$6�(F�.�a+�68q����:�:���3��P��4M7Vt �9�l�(Ř�p�������f����X�R%u_�UZ#�'M<��fа�����C~���W-�g6�f���n�Dd�|�[��4�Z�La|0P����]^H(BB�~�����n�QD���� �Xk8<�J�`Hw#_��=���;� �k�=���'gǥ�_�>[���6dU�bK����?A~�_#�B&�v���|�h��t�q��8+��d3�P�����.o����&h�FΖ�u'���!d`/ۙu`��w��w�A�kmz�dK�����]E�P�!��2�4��FG���{��/����G�	{�{����7��ި��B�p3,]Pu�Ѧ�y����ty�+�2��bC�f� �Q: 7�����������t/n+�S3E��x�dd3��
�<��*�9�^CK,x�Z��� �T7�kc~k�cyC��
��N~��0.�Y#7�eV#X�<ߪC�b���:y?��� ������$�J��wH`g�$=��gJ�p����ZHC윧�����f9�g��"�f]*7?Ǆ �ڹ�f���*�Ҵ�<���Ȧ?�
� _�����F]�9T0Tɍ��ӱ��s��A'G)gҌN����#�cڡ�[�i���>�x��b	K�/�ՙ����O�O`~$���uzzg�Ŏ8Ŭ(��E~���5��S�k<�[R��U�ԯ�.�u�,7�=]��`�.�3>��h;t�煵�]m�f5|�#J*m������,�ڶu�L�~R9��<7Y@.��v�x�RY��π>��8Uk���s9CP(�$��z��!5>��x�x�D���	�YO:76� ����@���d_ �5$W��]O?߸?p0��LӼ\�B����� ���@�k�&��V͔r�^:g�"�)���M)�D�Ck��e0p(]�uaAiv�$�U�Z9�~:�9���5D�I0��0���w�5��6T��37�9�<�Ԓ��� ��}篖���n�-�UW�9��*��U<,�c�_�Xj�G�Z���xg�"���
�Wz�U�|$���O'j5�.]�,�D��=��J6�V/�=����/7g��כ�	������u�$�لF����/�KL�@�U�T�h��m9�������C&��].������������gkƛ��	���d;JZ��hg�N�V���J4�g%��Y,տ bȤ��wΧ��sG5�*�M܆��t�	�ζ6s̹m��Jʋ���=!�}w2�w���>��5��kX�{I2�?o�H�b:�Wi."�S��ݞ�����:NZ��U�~y>�䯇�/��0��80����j��4"�)�I����4	\��j�d�~)�K��	��h2��Z�P�R�j���'s����j��+x�Ñ����g@���K���CN���N�BSvıZ�%F�/W�y[���-�.���/��.9	[��W{�0�P�^6f�jgc�!��7]-ŧ�.;W/\��0�Uul�3G���E2/�5���Dػ�M���Ʋz�ڸqgg��W��V�TU~*Vm��0��:-�\���U㑝��齍h�X3U����ޤi�u�5�ӎiC�������
	�\Sz�@���}yc-�iʟNzS�J���wa�5 p�wYZx��j5Z�a���Q�7�����E[�@��UZ�ŪW���E�R\llZ�2x��wc�;�4���=���0;7ņ�5xʠ�|SI��Vf���PMU�
��N�,p/9*-��3cx������Ԝg��U!S�>��Ʈb��"xcAi��u��Ia������%�������1i̙Ֆ�Y��k-����~�6��[?����V��W~�m�k5;x4q��91��ڟ��,��&:CM._Yhp/ jJ�9���fe+�RBS�����m���F�|U\�wM�5�U��W��H�G�+<�$y"8�5o)��@2�B�oC�qޱ�a��"����6�L�;8�xN b7�Ҵ������!]�d���I�O��`m���j#����+7�L��ʹ��#�`y��O0yx�?Z��0��4PG���:#&�aI8
��\(6�	ǹ����Qf5@׊�tb(��
c�!��H��y� 9�>(��~Ns'�ȑ�4��\�����ޮU�jw�U#���q|�i=Mnw�����n��
�}G}=&�0���	�-O�$�ҫ��<b��\���	��p�%c�����U�	�ȹ1��+�eBb���*>�D�l�sCe}�F��L�'�*!��l�f�J��*״Q��Lhyx
��~�F��;��"��գ�:���"��p�FB��~�,�IM�~z�Q52jo��0ڮ�9)j��Qj�
~.0LV����%�_<��}A�4��(V?�XL���\`�H������,�a�Y��E�',�JΝ�>�ZT��Z=�����ܹ?��~�
��ښ�*l,�Z�S��$t'kkڰ�-�����|��2Q&d�3�`A回�oX�I�� ]��{N]&cWN6�o���R�֯�4���!~��Æ�%��\�ň���Kf����uz�"z���1���qv��(lM�����-��s����Zs�@0���O�3���#����q�����/	���¨�P-K��ԩ����!`?R�)�v�([0W�Fr+�lB��Zr]�f���9�^F�h�Ht������`�N?�d�>�OJ�(������v��e�܅�rN�px��!Pu}�'=2K50O����б~:���,/�W�8s�,p%��P]P]T&�ko羺�[β�z��3���		����N�[M!+�'�1r\�
%h�U�y��+5 n6(|�z��z|MA�� ��F�lP���T�Tj��C'�a�g��BQ4���0���{#%eU0:%��.�SX��gN�1A���c:�J,0���eȢG��Ƥ�ϣ�r�*;�j�w���8p�V̈�Ɯ��x�D2��_|��#5� /���{�Z�*��(��Q��GB>4��FH���x��F2�ȭ4ӯ���8?���_���VG#�`�:�X�v�Ǚ���u�C��ҁΔ��HϹ�EKtҷ���a�X��,N�W�=�b �5o��]�O��ctU��u�;P{��W>��r*q)dq�}f���W痖��	�v
�y�[=��8���s7h�l�TD:Ur��4hi�&�o��	l���o܋	X�4Z�=�X��_p)d?S��A�!U�s���ۑX;6(J�߿�.�����'}�1��m��� L�L��8T]������{[c,ǎ���Y�����b%�P��x[��&7(�c ���~��N(�=�f"����/���崉�a\l�|�Y�B:/#�T%��/�%u�`Gҍ��a����Y��d�L�U@'+#X?=0Yꄩz�*���[�a��$#�����;�{�	�����VH��@����B\A���,���"�@�.t��Aqj���i?�(D�X�)I�*~�-E�^��)o�`��fF�Zi�0¯���8�{?ȣ�7����'i1KY�F~"yܘT������5�ZM�T�vwB��zuP��e"7�1�����o=����gH ��xX��'_3}��Rߎ´n�1��\}7|2�?Đ�-��x��T�m���Y�3i�߂�K&�A�}fĹ\1P�-�L5�uE�4&�/�Q��M@��OR����/w�T�:��Y�b<Ⱦ�7(��<�rn�F_��=��������Hr�!ٶ˲b��?���B��G�ֲ�u0"�[�}&�P6�\L$��0��ҝ�`ʷ=ύnQ��e߹\�V
���I��:cצsb}�b'�FU��U�J������1=D0l�'[��Bե��'y����<&7��/no�kRQ:�6xq[d��'�����^�Gc��������k��N�~l�m@� ����'�S����᯺Y=��q���[�hq�8m����f+@���V�ί�4Q������W3�e܌���s)>�����ݴ���(M�KT(��3��H���ǂ�?[I��h�ϝ'ZS�Y��[�T�s��/W�:��S�;rj5�}O&� 
��R�U`�Ah��A��u~���$d�(�J��rg>���j^����>uP9Ҹ��a'6]����� g֏��u�Hp���VO���Ûo��f���ǁXu�����i{r�K+j::6���T�e	�Wc#���i.ŇBR��&>yTD+���o�5'[�5k�s	����J�3(nem[С��i�Y��=I�ؓ�˼'�'�r�צ���jL`��R4`�|�ljhl��cܯtE���Ns!�#���,�� ���Yr����XE-�kж@f�;�/O��!�%Pj��dJi4B�+)�8^#be��+�P~f��w6��L>�s�(��7�Q�8(t�`�uUy�S� $AI��K!*�xxpgFH!��-e K�7�&U����TMλ��~��u'��<s�@_)�؇�����=�ڻ���"��c����EzL�l&�pQ��4�q��(E{�$&�..�4���D�/���̛Ʊ�,�8��s'.;oD�J��Zf��1��4̳����f�ה~��f�;��۰�0)��ԥ�=��`�4�!�_��b>���m(��`�h���#4��^7��(�����*EBh��,n���9+��Gi�գR�G�ft�c�Y���B5+eX>���H({�q�ЉxJ�M�Gpgu<s�"#�t50
'��FboyK�uL]x�Í"}�	��h2�T�4�_�j��;�T|�������\����A��em����V�*N���(�^����t����'29W��W�=��a�.r��!L�NHo�X)���Q;םu�m0�g��>D���F�.��bȲL����m��?t�$�
X	>+yU�/|���:��?�4'��Z��>b��n�QΛ~�h�a77q��*������3 2�oY^	4��2Μ�`���:�p�[�r>�H�>�S�B�ҿ7��e��#�Q)}g��g.c��'�j.ts�.|*��"Q�W�Oj�<�z�L��jG�v(#("\M�KR2����b��]����-��O�1,��{��3@ۤZ��tW�x�<��Ta9m����_Y��e.V�:�+��.�>c�;x�P�G��B����k�G ���#����E��2��T��� ��뜂n�/A�M�l��u1��K�BGO�N�!��cT�!�?�`���H<L��*���.���X�0��AtTh�ǹV��"��:�.>�m|���1��)�4���'�Q#)��M�jԯ���h����,>��\ïu���Όx�#W����^�pO%I�s	%r9C.�Q��y��`$]�ޱ�As�*����g�v~�d%���U~��c���2�e\�l	������I��C�0�>0��hs6�v���� .���r\��;̴(���B��f[�"���2�,�"[Gk�v�ds����ձ�l��UǗdL3�W:Q���'mC�>D��M�����А���J�b��Lж;��l�+��!�,�#�-��E�q�z����%����up�8[����Q��unq���H�&�"��.���Z��;�0�{X��;z�;�^c=?��m��[�-�?b��
mW���El|���@H6��ӂ}|�o@�5+C�A��QL��5��B��*���_o{o�͐;�
�i��!љ\��M�&���g�=��aQ�}2q���pv�<���W�g��X=WI�$�g�*����8R��EN����;��c[�CH�H�Z�E�ڂZp�M��lC���	�Ѭ0����J���Y�?�22"1���#�OZ�K�>ofLk���.�]XC#V@'�_cnjf�+�2zjCe�m��t�&�-\�T�����E�Z�ulw�,�u���]�7��F�Ӈw�x�_���m�����r�LA.䓀J�o���kMi��^K�b�W�#�>vR �'-T]�O�Q�Ym�{��Ƃ���c"[-u2YYO�T��o1~òY�Ӯ�����~1<���(�/��Lȁ�=���(��ٳ#�GW�,�(�`��Y�I`v��{-��i��{.ߖ삚g�Iry��W£ɂ�q�Q�~l�4j����V��E .���z�yʷ}��S8��bVG�x���aL�Ƿ}FV��}mֵg����V?����0'O	�iZ�၃X�v�D�������Ԩ�':��K���O��.le?���s��^[��H`n�7�E�c ��*�Y�ְ�+��E��8��)%�)�1�/ޯ3��:U���H��L`ء �MҸ�X��k�II�u�5wޚa�q=hC!�m{��f�7���h�T��CO���L�����9��g��������Q�D]��и��ex������PQV8T,�w�0_+�v���m7��)��[�sD��8��ü�M��G� �bYZd֥}��b��X�tPYl@@�������╉c�-�D�u�+��J\����_O\{�8�����*��Q\lz'ϓ�0�&���0���R.|DW���t�X6�����\Z(�2�ܡ"�겁|=��f?n�$-��7���[�<��-�J���*��e�Po����w]��_�]��M�sM��;(��;=��쫄O��ݨ���z̙�z��-��7�d����O)� ��-vw���\S��z�sԇT�%�_'�C#1��Ď>��J�k��n]��e���j�K�<����Ps���t�[S���A��bW6u���F�fyx�q�R�6fI_i��kl ����w����^��_ߎ��7"G�t�t�Y�^���ml��iX
Wy+�B S��t�iTH��t.�J�tŞx)�V����[�u���Hi��qY�\�K���)�'�b�'T��o.6��~v�L���y����_��-�0 ��ǐ�Ǽ� ���L�&�R���0M�F�{0��7�R�pS�s�O5�;Q�A(a�	�u1D���FE9�0�r4P	� �K �����K��Q��D��T�������b�M�Ni$��s_��x[.���ia�=h~�����ʫE�,�±�!��M=�Y���X�]S]0��}H�O�?`�w�^��|3a" �Yz����3q����$!��֑e�n�j���(�y,�ӊ�4�6ҳԤ��/E�4U;ȣ���q������w�������w_�W�*����h��|J�԰��.}����Uj�R���o_�v��Qpۭ���9�bK����(��y3n(Hn� �o� ��ts)H٧�t����g'k����V��سr�gמ��{�v�O4��:*�`乜����`cT3ц#
<�s��,p��Y(�w�J�82�3?�+��~nmd�H�a�1�.�w�"7
��_�Y�Is�Q ��R�J�i�U:����L5�^{��R�x�
�������;��W��Q5l�]n�쪯��B��&�af*u4˃W^H��	����h�"�ԾD� Óc�H�_u�UXY�<ʝ�x�8��v'b�޾T����z�%W��!�I�֠�]g����Q��7.fqn����.��㷄�Jȇ��d?�Ȳ	M�Ȋd��������$��r�?����9[J�t�y���!��8�%���_�;`s]^ ��됛�.Ł��E+�AmvY�pg<��N>��ڡ��l֮�C�(|8�[��Y#Sew �I��Ȏ�&_��fo2b7sO���1t�Z����c?�V�*p�nè���n��*�F�8%�P��=��-��o������'���5�IHw�-y�
(;<*&xj�WDD�sj=J��YiE���G�NDpc/:�X"��Н�MAM�G`ݿ�����f琡��\M�xx����fCd�:�J��,4�1��8�2�H�����{%C�HM \�Ťr�8/����D�*w˗���N�,���=Q5�� �H���ej�#d�Hl���vD�xڿ��ӝ�g�I�	$�(^��&��_���g�i:�ܭ���D�����*ǚ,�*8 �$�	#=`L^��vN	���:�z��fGX(Y>��%7i3'gp킋��)l6�:���%E��&�]	.�\�p?��(����@�Y�͕nĻ������5����6P��s�N8ow�z�}M�vM6��U�	��7:���#y_�W�~�w1S�V��{Aб�.�9�
�ck|>�]����m����Ub&C��p�RG��`�Q�����Ъ���td��a�cޖ�x��v�Y9i�9�GM5�Y��aL<�{����5�$�7��o���	��F�P8�/&�C�z�~7�?�ƥ�pOt�C���,L���8D�E)I񳕟������Z��b?�d9��p�IR+���jjN�h�
��[#Q�U&�����/��`��YM
;rꎸ=7i�AM���N�z�Io�o!�ټ.���yH!U�ja��7���+8��9��Q9ƖB�I0;a�{0z�
�D�ݡr�7�MTR1��@��U�|(�i�d�E�;�=e��`g0=w��g�����΢�fY�&�cXCC����/����07������s$,o�-ͳ��7���2��q ���.ǅ���g�M��tRVp�SܥE!66w���o�Ĩt�i���%ɀ?��+�����X����H�������A�z (��Na@���)��h�q�E�=Y@qua˪���LZ��h��]�����k�:���
'K%�<aE��ѱ��"%:d&z��)KW�}&�{���Tq�&��OU#�oN�{�� E�'�-o���MP.��,)VAvz+��@ì9ˠ�p���ɛ������2o`QM{k���h&���������Vl=ۻЪ�0�a�1���>݋�z�1��$j���
`�#���������� ���$M)B���C􃳶ց�D�J��YC�o��E �)((�7Y��"d2�O7���� q�R�(:lZHt�p׀"�F�AnESŶXI�΁B��� }���5'Dc�/5-��v�j�Qf�(.w���:Zs`j}c9=�^��5��
�)z��8x��0p�iSv�wn��
!R�eP�x�ǡ����::�{b��H�g�	�Tkt�r��8�)��M*g~���b���7޳{D��	v\�g�c��7jov"���8-�z�r��'M���I7�t����#��~��klĸ�f�����WTߤ�C�Ǜp4�H�������/��
�e�_���/���a����DIZ��ߊw���Sf٦�/6k_O��LVuNݧ{���ud�׈�mcf������t���kr��ʜ�:�������gE0H�v����+��l��y��N�Hy@<�Z�{T��t�p1F�x��6fV�G��6���X�1���M- fJ�& ������d�IF��]V��ttgh҃�\�x��] �|�v��L���[���L�+��j�hvn����@q 2���l�	��+�{��E4θ�rN����xDdq���������6 �!�`TYrHi�J/	�)�f��yq��#��WA��Xi=P�.�q$#�Oe��a�n��0��6ZFw�ǯ(��E+�&ٴ����yLH�Hu��&nZ�CWv@Ǒ�4��G��|g�T� �/<�_#�� ���ǑnT�4�Ҽ�M�TW\g\Q�{Ce&�͈��J&����P,�-���/�6��b>�q���#�7��XQ�px�����P�a�~�=?��>s��T�S���rE�	��7`2��D�8E����ߎG�U�y�*3Ǖ�P���_����E��q$A�FUЭ����)���7�=2��gͬ���n�+�f���BS�5fiu�d�`z��Q.q�\�;����`]{�!�ɳUL���>��p���?3A�A�li� ��m�jM���F��_�_�(�x"~U4�j�Y@~��Ξ�j��b��Uݿ݋�CeO�t	�����RO��H5�5#��7�}z��!���P!e�a?%X���`HS;8n�J�dk�yN�,�h�Vpq���/�)=~5�]�%CHH^�֭�7�f���F.]�W��\����+~:Sq��㯴�)�("�z!&w�ݕ}Lr��k:,d�L-�U::@�"�By~�f �Jٽ&u�Kʑ� ���i��ݘy�Z�PeEjJ�A1.rر���ޒ�X��]��h���o��~S<^X�0�+��Hp]Zx����<�б�����0�x��ӾͥT�U�A�ZmP�$8)�	�:���\^���p����Id�%�� GନM~��a.�	m��O�ZG���bkD�
�;���}ى�,J����?�����=X����K.mJ�a�H1�����Yxꏕ_��`�����Jf=�襩V�L�nH
.�~Ds�E���� �ψ�L��ǯ�����2M7w��Wl��wz�e?pk����l�kr�U3����6Y[���+9�,^E�G�"^� 2�;�YPwOE^tz;�tS=ek
z,�3��V�j���gzk�9r�bJc/�XV�7M�hc�
�7�k��9�E����?-���?!d,ĮFy�Iǋ�m�ݕyQ�u�����98��O�[(�֤������ l��TrW+NL$����p�ﬕ� �����x�Vvt��r^���v9��'���Ŏ_���U� 4rxy�+<<9�3wsꟕ`4����m\@do��g��6�)�3[��	���̠�OH��	��.���#��$^�_`���/���%�E�uUn�S�L�P'E83�9���'ۘ싕�/ч><Ũj��WlG[�C�����C�,A O�p��r�R�Å��#R�^���dBX�U�օ�p�����:��+��Kjz�B5�ݏ�kY�}��&���~�3�B��Q�+��(>��}����\GE�Um��CتwU�8j���p�#|�������2,�L��54��UVA��d��T��݄�)�T/2N����JF��[���ך�W�^l��zj#�s1/����\o��lu�kO�\�h�k�;r!��o��X�t֎�t�;U{?��i�j8H�l��4�U|���Yы��;ObX(�ԛϫ�y�Ԕ45�#�C�ߨ)H�6�x{��్�����A��8��D�#����I �r�*��~|�ʱm9����٨�� ů��W������h��^��Bp�2��n�L�xӛF�Ԭ�ýY��*�ƔfMd-^\_ێoI�Ʉ'4�6�IPs7�Ɖը�m��׌_C]_�G��ο��P`�<��,�����o$�]B3a
{���{[��zo������;	$>?0"kwZ��;1���j��UX��#�
Kz�4z�M�y�0�>���8��Nrآ��	��^ӥݶ�#���Q�ѥ�EH��>F��T�n�����,�}���:Js(9�(Ƈ��T���I�c�'��1h�-�P�Enq��{z����dbΫa����tˡ���"�r-��ɜA`FFܸ�\ِ�*�S�R T�=���sC�O�6����izvd�-�P2�q�/E�p|����v|��Dj.{�/�}�F�!ŀ�|����4�cJ��w��C�c��sw��L�n0ZA�5��)D�y!�y-��׻"��e4�l�.�N(
�FO�F��>%&v�|��JQN�zh�}u,���J0s��o���j�Dw��n�E���U�,�������c�����e?f�f:Mk��?���2�Ғ�T��~��ҧ1�����2�����葅?I����Sk/�*b�1z�S�aۧ��TJ|�l���5E�Js(N�a���x���*8a6	>�w��D���ب�`�9�;u�l��ŜNGQ�8*�;�,V�Fc���Ѭ^iJp�OB�����0$����5��鯰5�Qm����V� ���k/p�|n��� Ua�R��KU�B���%�M#�R��y#,��ա���ܳ����Z���������߂�;��T��L�8�/�KFVPV琍Vˮv�u>4Ƒ������DK��( ���m��_�]q������I��˰��.�E~�*rbg|��ݺ��@A��[��������L܅�yM2�aWG���� A�OT�1�Io3�&
�6��f�� ���A��gЉ�p�[g��}�,Y�d\�L�a�~Y��WK�V1zT�r [v��G�^�L��Q�Բ����1LpGiڃ��h� �?Jާ��L���י�}0��6]��*�c\��;a>�"�rZ�?� xd%P-04�;�b�\���g�A�X��͆��4�5�!׽��O�x�u�B��+Tj��m{!��Jۢ�F�<��NJD����V�D��4=�/(�[g��R��l$���)`�P��
ր5��t�<8H	O h}p{\� ��Is�� �*�]��<�]H�ސv��xV1�WA�B��o��t��y'�49��N�G�3Dz lW\��-������|]H�o�D�i�������.o{������k���U�5�"���?t~L'1<�g�iE�u@�8E`r����/�U��`-x-����K3ј �;j�G�Ge*f����>��Z_����DF0��\��#���U�A$�� ����u��>�`X
�ݣɂ�����9U^>4Y�e�vENz8E��H�ĄP��c�r4�ZU��|я��>|�������(��3#Gb@�'���qv�c#�����E�.�?�DV_}�g�����)h@��0I(��T-�닗n�����/7��X{�t�+.���,Y!A@�Q3�?&��Nb��%r��C7䍸] 8�`��#"%=k�T�*�:�RP�3�Ɯ�9�f|�N�Ȕ@�K(x��宷�FH2�D��_��Ã�=^���=K~����z��RQ��!yL�P/��'º�@k/��kI��l���ufE5q$e������)�Nt�l�����%@7
C���D�#�q�름����e��0X`27��] ����n�%�;��ȵ��EO�I��f�(�I&������/�ʲp���>"�baW�^�L17��lUd�+�I���UZ8ӶF��Ede
��Qf�t�&_6ڡ��3L�.�T��M�U��	���ED�S��W��\ۅ�.�df݌l�a��Q�L�!Df���p'��/@}�&���g.H���	�_לۈ ]�Jg��t��e# ��o�lH<u$��2�v�H<'%��h���^�̔�u�������\ǜ��~XÎ�z�F^*����L9t�����0�\�O��Y�^�n@��jyG�s�*�9l�.����<��L+�6jx.:�|y�¡��yqp	�E��w�Q��< �k��L��!j����FRП�m�2z��S��N&��}H��a��������A�r��̡T���z��s���[ۘ1�A�'[n�]���(������
��ң���	�l"2���5�<����,�QI��Z��a}T=��`�#k����B�@ݝ0ܟ�;1M��e��K�d��	$�*v���#y(�$�E���C���h��!�$Ӷ�?��f?+�Z�O�D��ZÓ<��� �>��{I0,ܧ×zj)-�b��*�"�
��q�)�sKuR���n����n����mf$D{v�zA��v��E9]��x-����_��gY�h72,�	���j��u%5%Z�x�xY���ca����fZ������$��Js>h�r���W�FY�+����9}�a3�I�YV�{��:�Coo���w#;\�>����^V#d
�y�S{�ŭ/M���c
R,]��Y�Q_�����y2�>�K/+���(�Ȗ+D�;5u.98��r+�������V�4���Ѹ���֍��#��xY �m��9]����˦��@���7�m(��X�YU���)<�J���N��b�͕v�_��)T�J�o����J؏�	C[�L�����4}�?"����h�8���	񊛹�yi���%^��D�{�p/��K�\��\t�ɲX��YΖ%[����t9 W���p���w��ܴ��I��2�S�w�����%/;Rà&��������7``a&��t��`�z/�	������*KGop欞�5r�����������w�_SElx���_n3YǁL�մyv�A�U���k���V�Y���p�~��U�u�GB��{ /+��!���>���1����=���Kuc\U,=$U`���U�r��p�pB�t�	�iz�&��.�K�:�:�L����P���n�qI���$�;p�����Q��c�E�~�����'y�J-1���:�I|ޙx�M�Үd�݈�z�ՍV�F�	�Z�4�
7��U\Tq�B��gn	�"0hc5C5ĭ���{�M�03՞J�:���Rv�������:q��JGȋ�u�?G#�x�PR����gp��_�hk�����hI�������fxոҞ�!J�ܿ�ϊ&�ܻ�m4d��"t�z�D	 �����v%���b9y�*[���oF�-����9�`�V�k�,mg�֎��Q������[�|r���N�kP��-�Uk�Gόg&XT=��SzV(�$6��@���w��mɌ�/�D����W�Ļ%���^�9	96
w-n�̄��`��ucV�ܾ���:�3p��;Y\�0j�$3.z�l����8�HAE{�M�#�ѶH,*��Cw�U-�)�Ea"��B�7�6�B�{�uW�Qپ~�8τ�)UX٭������3��®RI�K�i�拇����z-��Z_ ��v��*�'1�|[ �ҌhZD� ����3s�y��(�V%���e�;n���n.'���i�џ��.�'�aG+z�ӊL0�eo3���zp��!9�;��E��$-�ƥ���0�b�PJpn�!Q�h'��1h�8����_+��JC�m-����<I[/�fU�,�h�{����\:!��/첈���a�$bO��[p@�����C{���#��r�����)�	B�������Φh���&�`�"��.��Ï%�f ֈq�燕4	�(i*}�%z�4>	����;1��5G5Ӹ'��>�D����(Ŏ5�*A]�7�O������-��.zUR��f��S�ۡ'��њ�X��
(����xF*!�em�/؆���z�s7yW�@�cR1=7	��_
����A���ͷe���}�D^�M��@&.ѕ����,����� ���Y�7��#½��_{_�_H�f���/���V�Fju#�NŚ�qV�̄���Zx1��}m�7��g�f�:[K3i�o;9���a��= �50���D�֝�>�M���v�Q&��64ӻ��}�����O�L�w�bF���>_ǫ���jq��a���T��d��L�S�.F�]�*��",ND���[��^vQl�??chůQ����'�$0�1Xc$C���͔�X��m�ơz�1�[��EGt�U?e��2��_�O4�!;�X����6�r��(Ն�5�ֱ+�#9UR��m��w%��#�����&�-E�i�r	M�*[ �ҡ���|�f]r�f��d�o)C��l��Nk4�,O_���ɽ��	�p��`���9��jn�5]8J8��%\�[�@G���SaI���V����5�S:�41)�TG󐩆%����#�	.�@�e��1}������م�Ɛ_���f��� C]���鴐H�kE� ���s��B�����9�(%�:�-��-��d1m�_�+$�l���� �z9���� 4K�������~껞��rM�����e}���~��8-?b����͔g�M����8V��>ߌ�~��i����Z��01����}���]*�t�a�{���j��Z���4/Ud�
�΀c>?�A��agZ�⠗�~e�R)g���f��8'�oA702��٧�aVV�0-�0����Q���� {v�b�Z������x"H�E�lKt�����n�!~���V��o.9FW��EOJ����/����w+`�Ry�ם����dHA�r�˕��W+�:pz��¸[��1*�Ou�x��:��n	������BՒ^�3$�Lt臦���*���T��W6:V�~:�3Y�m&�W���H�2��BI)ճ�]h�t�N0�Gޠ������=�~�}���d�"���i�)2c��h�W�n�G���3f���$���n�8�*�<�l����qkI���E�������Q��iFcN]��-���>�Y_.ܕϷv2Ԗ�ch�|q����6�/����I��m��S���iC��3�̵�գˤYg�+TIo��
<��<Ǘ��eah���e"P	�M_�K���@*]�(L��q�C����Vљ��j28��m�3��+�<�&?�1(l(R-/�[XO�#� �@w��hVh*M��bdq7��0�g�/�Zb�T9������7���B�*�Y\-:���@8ɇj�jM�h�Z��je��}�HΗ��b�M��Z��(X�ŷf_#r�7ѿ����0W�C+j;�#��Y��MN���|���ox���lZ����.0O2�mx�@4L�,������1����y����0?g%܆��{7���u�	j�*\����%L�T�粊�xN�d�^O��xa��i�P�L�o����D#g5;n�)�#����<',R2%l\
���'���! j@�b:ɹ���=�/���VT�Gn��nQ1T�(�>��Q�-�1;�@'k�qz�����X�{ݭ���$��c�w#�T��L94q>ʼm�� �,��S����'�9�bY�ъ�@�>�u�o��2��|���b����aq�}��n'}S娙��qK�"�����ɦ{L1�}�'8� �֒,;�g0�!J��t����p�^����˻B�r@���ʶςoq2�K��[��lؓ�#�
F�L3�[c�],+g��UtL�^N���m�j'kN�f]�K����������?��8cs�TylԾ8���c�Ц����䩴|��4�6Z7��6����9��Ñ�G�M��N��ퟴ���eEz ��ܓh)��v�u>Ne��AVClX!�q��H��b� g��&
�q�
� !c��+mj���Ah8Y�aa����
G�b�(����D��[���]fq��ē�U���G�T$�����ηl�U-}�9�y�W&NX\]�o�6.�4-�KqPH���
��E�I���L��>���g�~�ir-���E�WrIz��V�̶9f�_/�0�*���M22W3�]{7u�$�f���Yn�P#����7J^�:�;�p 5��4�T����q��T�ĲJb�g�	'MVX�D�댔.��)����P���v��E�P!�4���"�G�o��kʯF�v�i��/H�ѫ�l�noI �|z�V���th�]v>5����l�ۢM�����>����%5 �z��="��@A+��O�ŵ4_�Bsݯ���x/�	�F�?��tS��'U��P��Ѩ5\@ER�x���G6�~qM.��}��@ʧ�
O�H����O�&��������qBؾ������q�Er�������^�\̕WfD���-�xWE�3:�P'���⛇�3���zi�͑T���EY�R=EMW�c�.ItOi���B;�����fw�&�	�,U�|M]
3���u�R��D�Z�A��7|@�ܯ�Ұ���.�`5���
$�x`�w_ۛ`ȗ�3i
��D`�Ty)��5��m����C�uV8��5-K�y�@x��e6&(�|��<Ƹ������/)%�����n�t��ǎt�{�4����{W����l' �/Y�-�:p2��T2��|
�a��`��o7FFD�<G��ks��y��1��p���%�ԧ�����-"�>r0��n"��u�Wl�tp�3�f���C�|�8��Q}%���SW^"�n�RfNҁ�׾�,���z�g�?���S��U����c
Lk���u%���C�O��c����K��Pt����D"�F6�-F��6���3���F�J�|�89'��MErmL'�(7�D3h�¶57a�،?0|�{���� qЋ����^��;�L�Zo`�K�&Gd�����$�E�L�t����#����`W\%��?n$��矋3솺��Ա���[�]��`�}Oۛ�f�p��'���_���7��S蓥\�+��Y{C���6�#���ba�V�a�:]u������8�Vg&�M8Q��Q�����s\8�#d��E}��}.y�A(r�/"1�4��?���[(� �D��������fd��NV�c�4Rb��n:,邯��
���l�gqj^��diY�,CY����I�F{gS�F�G˘YZm4�QƀA���,�!Ȯv�;KM����-�FQN�����癈�5�mE�x�i��R���k��*��/"4�4a���Q%d�E2ǥMã��~�J�H�7�2�$���T�~~�bӈD��/�갚���80�BhC[0��Z9�X��r��r�=��ز��}(%�(��N����N��E��=�Op|�7\O�d)��qa}̛7�)�����~3�.�f�o��(D�),͟��B@ ��'���0%-dy���L�b���EJZ��]ځo�"��Uj�"��o!�[<%&��2�@_�ކo��:�ﭐ����J&졠�6:T�𼘾�\&�+��ʁ�f��s�����,��L\��1��� 'zO�&N���o��z�qFQXAV�=�e~��r�E`k��<U�ǠP|��Q��aK(�W�G� X%a%�<�Id��uw�Jk���'��kg���)�-�H�Y��g����m��1�$��#~��y4�j�$�_����rDe�D�J>����p+������L��k7R:\��-A ڟ�в��Ҵ�6G��X<>�;U7��f;�Ua�} �sd��MU�Ǳ톲j ��[6�#�N����W��C�F)x���n��"�I��J�?�0;vN:��,+n��-��C
;F��|���׾�����Q⼟k�[�	&�R�{H�#�A]�9��7�|8����!-�l���9> 
�pM5f���r��"��3-���ƶ Y<���:Mp���R�vHpN��VyŇ�5HZ��,�'8��2�(\4���y�$p}�N#�`\+�ٍ& ��T����\H�h���'�]���ݡ�w���[������Y!�K<�}�-��`����
N�cE��ًp�H見�2ؐ5/����Q�&E�.�J�f��&	
����T4���dT݊r��5�s>j�'M݇d���x�hZ7{�T�r��<�dTM�4�z�ǆl��1�S4D��!O��%�j}�����14�ڥ���Mj�5���*W6����9˫�?�&��H7���4���ɾC�(��jP�Vf>��Ut��Fʼku��j��/�?��'�1�|���M������Ԅ���Q�{��g��o	?��\�[W�^e�����@�C��=�p�J��ix@]���X�Y���qc���!��(b؜^��r���Q5t|���9������*�T�r7N���.���sX\m`�x驹�j�0fO��S�����E._r=W���n�X��&�R�(A_��f�����t��jմ�[fiS�����;a�}����?�)�a�zR�9���sE�['�TӎD)1�XI1uvq�OuZ ���O_�dϦ�U���;�44����?�� Z�f>����(��67���h%��.z:9�E�5�/즸����TuOr;����o/�����.� s���S1��B�#�)��nB�q��n�c���a�����2œ�Ĭ%'�H�PY-\�FQ,w��:��/�R��J���"�v���q~�Q5�>9�2��*���(����6�Ӡ��A�<+����9�/m�8���3	Cg��o��6׎�t}���:�}�K���~K��ۼdzPb��j#��� �g|(�<s�m��+���]�����]�̩����@c��nq���O�
%)k��p��KvA���Ψi���\���f��;�Sg���b��O
���Nc3���l��΀��ǽ�\�eML	�NYU�+}�&���}vp&i���H����u�1]��l>�P��v�S�a�.״��Mk@j�=0�����C8�Ɵ�w@e���յU@H�D��2�eH��;���g>�!ⶬ0���W��NE�g���$��6	�������Yuo�#��qw����x���#$�;�
��w�s�D��h՛品����y��f�,	�/�@� �"��'ȫ��`l�ԫX��'G��Ol�j���R��Q�y��d�J�k�f������ig�1��\=r�}+!����_�)L�@(b
yye�	w��G߂D���3eg	va�`O�D�y���:���+Qe��S��7���1�q�"�1z:�*]�����נ��]k����U6&}�.Yo���j��h:�����'�(�g3���e7�pt�v�Ӣ$"(��X��%��b܅�G�b��[�������8F�Ǐ]:�˼�r�-0���c�r�(�ai�(�E���W�%�o���0(Nݿ[�L���C/Bn�-���}�����G(�����տ���o�8·0Ś �ƹܑ�`��� Q���� oaP2������4�,��M���f�vW܏
L�C?�1K�q�P���"�ʩ��=8�#躍�)zE�n��&Ш���G�azL*P��@M6o)ۣb:�%����c��<�|��sq���~����88��mp�hp6���|��3�0�L�4�n�,#%V��6�s��3��D����j� o������s�Ʊ/��:�h���0&7>��8�z�Ie��{%�RQq����DT��u�cm�z��/7U}��k҆KY���������X��nL��d��JO$6�@�K�TʓP�X�qA�ui����;/,R��p'��һ��E��y͝��=�ym�`�܅V���EӤ�|�#���t����e5�t �w�EMVg�*�c���<�˳Z�#'h���\�qU��(坆E��e�m�w��3蝕��{���dv�[!�lq�w�fc+2S���m}��r�YS���{�(C]����t��kV4x�K
v�4#s��u}�VƆ��X���Z�]�w���oK�QA�!m�T��i�&�r�ND�������l��"H�=��#��P(ES���V�3��n9���s6^Ebg4ym��7<|<�5d�9�~qHPO1?|wJ�)��[L�U1��u9���eΡ87��H@���[D딖6V6L���$�2���'���0�E���3�[��m������i;� O�1�=�p�b[B�}�.ܥή���Av�4�e}>��!���j�����Li2�h�8,��VAa��P�i��)�X0�˲����j�HH��Ϫ1���6�z���~��:���lA��A�ل��c�7���b��&���I���л��N����<�ϟ���E��X0�AQ_CH�v��������]�Z�2��oJ�HQx����A[�#����e�D	mU?ŕ=���ϋ�+��գ���v�" �������ީ��[�8�@�|钳]'�Mt�1�`5n�P��:=�K�����z�����΂���	�ߧ��#Qt�1���ڷ�zo��4z�\:���a����S�,r�z5x�o�`z3�����J�)'�\� �䇇t��^��;w���;Kf�An�6�s��F���x�5�J��� <��=���r*��6���9O������ �8d���� Ad��\��3���7���?�sI�L^�`����Tkks~�Y����]�Ee���n�=5�,ɣǃ�q\K���V��OM��$R�U��F%��)�����(3@���?q�9a|��݈���p�dh���b�<��)J;�H8��5/�i@@v������)�U9�ud ӂ��!9I��i?�R�%�4	1Vq�\�Ա�y�x�',l֘OŤ����sPu8~��M(7�!Q����� z���u$<g�.2�����lM�	A��N��ڲǳD�<i���/rn�O٨qEE2x����aX�������0ؤ���
x!�\��Yل�>eT9�z��m4���m�_R����{����?V���Y�SlQ�U8C�*e�<!Ja �I�m��V�������	��{�9jK�����g������QoQ���z��x sa���BV(@K��f��p=0iN���\��+�-l�'��o%��Q|
�}�.�G�üTYމ>#D���wY��/!-su-BuN��B��3]� �X�י�,{Ց~tZ#�8N��0gAf��Yd�=Jky��
�BkI"���5�Ǉ�u���5PJ��6���A��*Dox|�}B�;�if��rR�X��-jMt���B�E4��:n����D�HWC�`UкJ�Rq�k��O.o�룂�qL�k�9�!�y�X��^s-s#��OouW\d�4��'F%{r3]>r�Q�2��� UِL�����q{) ���k��ŕ�X��!�p�r:�(U+���׮p�ӽ��%��,�	����B��u'z�3R����v$Y�ν_��(ݏ�;�=��jm�ň&��g׈��n�ĵح�U��/�a8g�H�q?s���n|1��粋�L��")b���bI(Ew�BL	j��uc�T\��? �Eqiw��&�wiu~F��f�a��ic����a�)0���H��W
�[!`'��U��LPh��w�k���~s�x��@�s�+V2◹���,��yfC÷�bV��F���U����5G�i,���䓖&d�'�I2�n�}��#
3��#���>^�ql�j�C�Q
س�.�0:V�vDu��O�CQ�S���8Z�Nu�C1���C� I��5r4�$�E�#C�ˎ@`ܡ��~FB[_L�	��J�3�0F��E�u�,��/uj�B����\��2����&͏����)��8lR�$Ǚ�q��I��c��Y��j�nq뺷�I�6�.,^.p��N�����'%��}U%��Jg�H�Pnk� mN��æ�>w����n�|���
�(�n-�ܛw�����! ��z�<_)F$�hѺ��-�Z�m_�m�oN��WFS°��(�a ��(�e�ıq�ȃEoS3qJl=���oئ�F�9(���oQ��dKK�c�esI�|�d �Js�
l�Ў�e��/�d��ֵ�����šp�>��c�|���	����qb5�^4����pǏ��Ql�Ժ4ӭTl��	j���?7Ҝ��7�ϊ��ϻ�%�V�ϷQ藬�S�������ח{�?���7����ʗ~�����m���@�1ɠTe����m�;�>��5���!:�l�l�4*�N'�$��p$0[�!iV (��0W�,�SD��y@Tk]\r��[�R���WH.1��@�@����8����Y��O�ꔥ���(xO�%�_�*��j��R��+Q���ͦF�
K�L�X[ѺHq���VƉ*q�emz�?a'�S(��w^�4F���q��,��q�&����x�����-qgƛ�����>!j�3�r�$Wr���e簭!���y�	w�J�gU�ny�����������x�^�i&ܓN����t?ji��v/J!�'���('���ok��5@����&_}"D�rw�V!����s������q �r����!
�ɀ���"�W"�a��0j�$4���1�P�`'��N�4�G=�L�M���Y�:��E��#�6�gVwkaK�7>���v�UQ �$�}���I��6"���+; [��j:�#�w�9E:��8G֖'��"�E�~�Ӆq�*z+ӻ��d�^_�2�������5�[��#i�j����} ��L	�8�u��)T�K+�g����p�g_%rЏ.9�v
$'�g��6�ሐ~3Ky�o��:��_�3�hD��`_��1��9�j�%8�:)���%�bb���'ksa����5�,%��3>�\
.4��HpW-�+�m�a�Sg�@dnޏ�CK����9��z%N� �}rQzx��Uv����?w�Hm��*Ǆ��
�+Җs�&���H��aR�n��%��p*z�#6S �O��W�,,���
�y����+&w�z���{�=�Dc�hkkq��slT�7]�O����N�3��|��'����ZqL�e�x7�4Λ�O��7I&��[�d+��Ek@1���P��R��������V�07�G��lV�u��q��3B��b)DZ&{5�pX�鲼_�Jd�7ss���%�җ�Y�.�΄(Œ�6�.�S.�~�_Y���;Z�@�m|�!�������IU'��1mʿ��\65�g�3G��fF,�wP'�����I@�q�-K�^'"d�44����H,����\
O�����X�gfP=�x�����We��`�[�^�V��m�ʞ�KC�=��Uu��]9��r���S؆��@�����L�a��՛L��&�s0Y��K]#:�h����o�m�5�0ڦ9�3&�ټ6tz�1ԍf�U ��`��*�/�I[���x�>�砄mu%�i�w�:�Oب��8첪Ӆ�M���Zm�Y�֩>}b�ZX�j�H�>r��5����dk��Jw)�P<vZi�7��)❍@F�\�G*c�(�Y3b��0 �E�H~]��.{W��>�V>>����ݖf=�#��x�a��2����M�ʟ+����l8�O��]���f���q�ᦊ�c�O�"x�	""5��ｷ.Y�Ӱ+j��n`��t��jp�������B"�<D3w"�3�H\������iKP�BTxț^������ki�����,E;�\�3�7'b��1�C0� �i(����K4�؟at�~ݖ�BS���5��w�`*ƫ�V	Z2�gT��zN# �y���8��1Zǟ�����$:ۭ�[Z�ji�|,��Z��o�� �;�V�$�
����*��,w�3��w@�tX�C����U�q5*� �H�$/��龮)6S�_�����2���O���Nj�a��8��I�3��#����Z��P�YT~���/�ps��t��x��;�V*�oX���}A\w�]R�8K�t�A�Z[�i�t�5�@�r/ۺ(�?=Ae�l�xY`X��N����M��w�ѐ�}�W�����E������tr� �ϯ}�zN�/������
;A�8J2t? $��1�܈M=�a�#79��t���LvBs(�:���VB 	�	z�.��8�!�a
P��A�g=+r���ôW]�>(�"s�h�J�O�� �=u��#�w���q�Rދ5�n;��au�h;g��Z�{=�u�)��7R�J�PF�)��ܑ*#���y���N*�N?��&�r�i�pl���e4Y��y7{�����&Ƈ>������:���K�_d�WK�9���/�:�7�PðD�KxN3�S�����Dw*��΀� -��+�����
L���B�F���=�~�ٌ���g��^�rBc�n���0�YoGm�U��s��Ս��﹇� ����U�^���ʎ+��k�K����2��l�2f ��F�0ܭ�,�� �8��0��_
����}Hf��G �`Q�&C��)k8V�է�èd/|��d���f�ɹ��YB��&E[?*���ˋ�ʻ�7��~8(��璳��K/d����)����"�� ��C��:k/w������x����Hs����1�À����@��O����F�bWh��A����|��8��j���J��4Lf��hrf�9���,�����4uD
a-#d�r{����4���-2��G�o,��'�����~<�1$[�v?���ѥ�8@����lO" 5N�XR�ã&�I֯G &�%��Wn����%�.mSU=uH#
�H�*S/���%�d��M*��ޗ�������\S1��=�d��Y��X�R��7���6kG�,�Q	twM}��(!���z7x8�y��3��E�y���t��Y�z�Ng��][ɬ��9�eMS����\�OW�PP0%߆�B��y�z8u��{S3y�;OQ��R��Ҝ���{J��~��K']�u���OLH?%u�)j� �C�w�2�X�`H��p��y����4�w�aL�A �_�9H������/���D��)b���n��,Lo4X����n�p���{|d������T~.�{(2� ����ZR/g��J�����G��:~�����y���Yw*`�g�R�
ND��������N� =���B�~��3Gl&/0\�`��U�tC����'J��f
���U�0G	��:��;��E��e��U��ʻ��OQv���M|���k��d�\��>��<Z����LPTe��㺄��͚�u<Jv�Bn�+ˢn�'e�"�@U��.4K�Ëh�|�G�,�[J�e4a�z}�A|b�l�N_�8�p�K*V�z�,a���IIA0b��_��T���$0���d�!�t��8l6����:sUS��ޢ�r�*���	���̆�6�Ak6�%�F���Y����ބ����=ܬ��`o��������z��H�:R6ច|/9V���Ǝ�����u���;Y0�-�	����Zw-�ȳ�J@��`�� �IP�R�D��1��_���֝}u�K�����U�)n8��p�V�y�?)ø��ж򕪺������C<�P�\g7X���{$�+��&H[7qOrh8�F�F�4�+Dn�������+\�,���!i�>AJ�Nv+h��P��z������ ꁐwΖ 1/���T��\ ?�ؙES��<��'��\�����P���ӱ�='B����#�J�\� ��F�o��O�֣��"����s��"�"/�I��w���6�*������[y=�S��:s�S���?�N�m�D�=%r��������Y��8��69��}���~������=�<of����$:5 ��@F�����/�$M%���1����<$���:q����?���J,���q����F��k�CM��ש���4I�c+@G'���j ���}R�vq�Z@yc�ߓm��jD%MQ�
)���̦9��{h(�$����xET*DD�u��*�=��wh�������Q3�S�4u����rp����cW��+����;GU�MW�ͩj��-�lQ�r� �g�}�ׇ�f��-*�N��#`܊��O�?�*��m�x���� ��A�s��M�wBZ-Q���n��ys� ���09��٣1k"$�GPճⷠ2��!�R`�P#��?-ODFY$������j�m%�h+�_�S�a_�s��&�����$�n�lՅl�Aa���ѭ^�,쁆��<�ZrIǼ�M��P�6C�(����iJ�L�[ҭ���g�R{i�o����_v�9Qڮ�FS~�D� �nF���\�_W��_tٰ_���`�)���%v��� ���Z�R�nY�n:�`�PV��'����hp�������lQ��ެ��� b��wa������p�����љ��'G�G��j FNO�>�j��_�����k����EܒA�!C��d���1u�w�ĺM�И���!��n�a/sFf�H�Ӯz��)[��Roh:��Ș�pࠖ])#F�M�pNך��{ip�98[6~��l�P��MH@���U��>�Ҹ������M�4`O��NG�\����✙Jd�nvw�:yH�c��F*�pc�(l-\|�y\WM'ȟe���4����)NQ�=o��Ԩ�u_d�v5/�;�����>e�ǥă�mo�A5.(�[����c�©��p41^�x�u�/^Y|����[�מ��	�O6����x+����_\N+l$�<Ӛ����S潡�R<��V:��(�ۦ��uK{���Fh����ŻJ[��6������o�+^����=�A�-��>J@�\-W��Ņ���}�3�c�=Uͽ�Tj�q?_�d�Tfߨ'��葱����Yf6��c精�5�9א7�/IQ�6�����?��N��5���R~>$���x�AῪ~	�BL�0g"��e��r�x?���5��:�f_�>�@s�QI����2�Ha����'"@6�,Z�a�{vEIbM�Q���Я����;�L��IcW�#h��疊X���g[B��s��#!W��S1�~��w2� �}�=�n{:��nE�/�	�h����irt�w<d��m�B�������Æb�n>��B9d�W�D��5O8��3�����8�������o�e���2ς8�f��۾:���Dk?Hl[�&��{5����er���ȅaw�01D�E�.ӒM���,���N}�J�����A����=a_� vߗ!��n��9QYC��7;v��{}��yb�V��X�|]�tb*z#���n��s����+"h��� t�^cxz�-&���ϗm� �D�e�c��'�iOp����Hm��罊����Ĵ���o�2w�ȱ�Nu�X� �����l�M��#?�WICX�"�H�,c�y�����Y��=?����� ��t�A\�q4Ϯ�h~��d�@����v��NE�`�
홵�SlԢ	��0���#Zw�w�P���+�b��'4�n;��r���<��Arx@�K}�K��Č)���{�ؠ�R�m�ԆL2�xr��^�N���p_���E"�c_E6�5+#y!x��%�6�B��;R��y�%	U��VQr(;�o��+A 8�2d=y ~1��Ӱ��bdv<�X��&B6�S�/�tK�������x~4��}�N�Yf����J�ԣC9��IX����K�[�e>髞�H�~ǟU����l��i���R�3����_���Mn>��J���(�ȷg�3��]N�_���'>UnA�z �;�5���M�vsP���Ƥ���[�@�R�������@m�/���V���p՗���'�_����hw};r�C�m�o��%vBç�� B��aˠ�7�P�|}'�x�����y���ҫ5}���B��N�#½����~���Q�Vp�Ia��=j�&�g[?���(���<��xԿ�iQ���6��L9n�*��BNPs��-83��_�0�1�����@���n%�Mkw%0�`u/�(��$�<P,�Y�z�%(܂M��F�y���	��P�W�ډ�mݑ�׾V�h� xϻ����#��� �^��:���+���\��̮��P�Nɔ\���xȼ��0�]�:7�h���E
���B��X�{x��H'f�wmq�8O=��&��~��*K���%iۆ�����R��*:Oݔ|�nN���FSr�c�O�7A�Y��Z(I\��=i���Z��\X�i�т�2���PȆBˏڠv����y�%;
:��[�����`yo�8P&�3'B�kU���36�s]M[�v�
I�uj��)�	A��$L��O-�O���h2e_����]���K���<kv81a�лg��E�̭�R����J�Z��"Y�N�<�&X1���<DHq!3������owi$4*ƥ��Xʧ`{��x2���
S&�D<sL���.��Kcp횭ugm]d�")+�H8V)�3U�؛� km���n%���Yg
����p#����	"�.%���D�Hձ�Bِ$�Ym.t�9���(�4
��3�G#�6���4���o�R�1���A)��*S0����V��V��PQY�P�<H���
 ��ֺ�D�n�-r�O�s8ښ_v�鈀�B�^"/��Bx@�Y�n��H�b?/��{-��Y&ӧ�8�Q�&5�V�w~B}q��K|)8�梞CEX��&�ͱf�c�͢@e�Z>]�*h�SF`��� ��nO7�,����Pdh�� Ĩ�`vVa��������x�����m;T�1��#O�Y)�A��	�OFS�*�Zv8�vE��7���?v	U�
Fⳁ��}�^	�a�J�F55����/.�d�
9�����{y{�~'ɯ�F�Y�)����Z�cs�Ս�:g���'B�FD�gS20/������ٝ����u\�U.j.��]'B�p�|���9�K��ݺv)���#�S��	n%dς8G����D������F��eJ?3�J�E�������K�F�nl�`Y��e�:ê�j&~�g���m<$V�]�9��f�����9��;X�+񩷞�3�"/�w g���7l��4��� 7Ʒ��.~�FU�9S|pMD�󖸩������M�[m˯ŠܼK�h�4�l�h�9wa@� d5Lr�i�UR��_��Ф׫Ƿ���j�v3{��F%7�o��T���'��w|�M�oJEnif�Nƶ���ū�$}����
�u�8 ]���`��Iw�U��0 ��*+��,sp�5Z�Ⱦu�y�/�v���H�Gm�TgA��O����l{9�w��	�R
,I��ȏú v�2�\:�bK=�[�����l����V���Qֿԃ^�Mq�b6�&���P<���ID||��Ô`�,�|``w���A�'-�÷Ω�W	�:�BY�#�I9�`%�W�S�.�.��|0���~B�;u���5z����P���6�Ϣ�0����3�c�ٖC�vySO�r��`eb$g��$�< 
��u^����U^
�A{�����l]R�K�Î�͖4��酷3����2���"b���	�+��;���>�
_K��/ޱ������d�F�{�e���"�B��ED�G�}z����sH�ޔ�.`D�1#�~�)A����5"�?�P��@gr�_��L��4��4���{�L5k��HV�Z�쾫}N�V�Ԭ0�C}��}��L~��(���ղ˓�/�t���N �<�q�!Qt�A�?
���ڝq��x��o"Ե�5 ��2�y���0���j궪�k_���@�;+�(�߬��e#'Ng?��Y�6��
�Ȭ�p��W���MhB�G��d�#��źv��4_ �$��q���#�
�Te SX��μQMA��|sHe��d� s�6`c�m�pH'��tK�Mش��}�󝘉��݇��=����׾GT�h�5�%b`Ya�^�G����� H�ܹ���w��u��]�r߬����71���zYO��wD틥�;��G{PbE$��T�>��_zQ��̧� ��CA^�9��!�5@�b�mo��,H������
�h�G��k����@�VVx�!���b@�B	 r�*iI�K��L���R�
�9���+H�鲵^i��������pϔJda�x�^��{��4�#r��)�>��ݘLA���2#�KJ(8>��K���
���!f��x��_f��5M`0ȾC��k>���,[.AI���F�TpYd������]�S��c�[�gn�{�V�Ы"E%r%��æw��׹y���y�f��CV��G�4u��?�멍Ĳ���?^a,�� ']�=��sk.*�A"�(���Ҭ��+xkp;�`��m�,�ʗ����ɴΎ����u1|z0�����7��	&W�%o��\��:�؟�1��8��륬����v�{1�D�����-�r�������ǩ���s�0}�"�U��;G���d��eل��+F�lr��`���D��Ek󓆳7m.�"b�c�{`�+	B�4l��#=]�4tq�QL��-,�{��踨h��iÌ/�uH�s
��nHY�-$j*'��tm����:3f}��BhP��'�������|w��N�`��<�#�@#1۸�b�S �8u�E����]�T��f�tI�O}!�9�0Zw:n�|BY�J�M�&�N����MlI�x֦�v�����5XOX��_8���x֥����@�|��?rp�����#�c�AM���c��y>�i�^���ٗ}��ׁ)}��^�iwJ��n�⟓F��J��0z�bl�&���%���Lϝo���7+B�C,�H	|ԛ�A�mb{o'��2[0cG��L6k��G������Ɠ��?2淄5o�ql|w�ζ�zw��改�}%�ȓ��d0��� {�qt�p�M�O��~یB����7v�Wt�E>�]o��r��-��򦄻��ą�F���>ԓ��&mP��(�u4!�Dq�GA�.�?���y%N#�B����ut��Y�Y�dV+�,c�x�*Xq;�D�_y$/Y()����"h�u(	[�"�I�-;nU�[����Q�����כ:Ok�LߧJCH�|axP���G𒙆1��&����$��^|q[��pw�ZZͨh:p��X��o�%�C�� �n�,$��œ:Ij����DT�m^n͛�w�EP�����k�FP4H��FcЖ�����
�H,q�R� ��c:!)�_�"uNpb[bή���F�]6]����u�:[kg�9�68��H�"�
K)�w|��3t�K�N�J��焩�J�O�?��D��p�B<q��	ˤ����K��>x���W�����>��RB��A��p�]��
���>���TY�o��ѧ����4����(��9�n4N���-��.��Vh���Wς���5��څ�(<A5};v Ax8�\�
�����l��6:�1��q��M�e$Ysi��5A.os�C��W��
�?����e��p���B�X�X<��WG���i�L1b�JfZ#�[�aj�T����bL�g +ᥱ���+o�߻ec�b�U6M��B׉å�Bj��&/���n{��ȗ���4�����/.���(j%J���4v��tK����3��M��f�a-x��VS���F�۱{�L��"��3�6!t*(��*Y\�ʮ�{�r�ԡt�e��Du/�I�*��Px��k���6�#&;�ᮇ����đ�h��#q��We��gL6Bn}ro4�@\,��1j��R"�,���u�Op՟ں�\U�EBS�u�<
��5Hx�o/kR��!��i�5ϰ,{��>tO�0@�bZ~K�v�'�29�U>��^}�:�{d	es��O���l�<b3!C����C�+tw74E	l`N�ԃ���b�����	j8����С��̯)�7�`n�;���i��n+պ�0be��H��a+b>���x�F��TH�ͥ�`�E�Z�R��L��j��1[�R9�*�,@�ȼ���$���:zG� ����1��2�4.g���?��h�����;�-5s�:o��!OW������mW��Q)��Ӑ-�$����F5�-E�Gs�M+bz6��'�Հ��E���pm�p�x9��������5_g�ծ��i ��� ��0� ���+�w�^��j�xL�4�ez��&�q�%��0�>��.j��11�b^)ҳ�9�'��nyB�"�:�jV�f��E���p��'ŗ��:������.��0�B���,Fg�`�`�l4�J�I���լ��ӳ=:���:V=s-��>���?&���9"���}�|nW��}��Dt7N�O��M(I�tC� ���, 2t}�����Q��+mo�8������GǦ����lʪ�M������E��8�9��ö���f	��&J�h������mtp�3<�8;���+��2\G��cӎ�E���w��F[%`�#Q���g�'����Uo��&l�0��zK��>�%�Ȟ�.�	�`�����IRiM�K˵r�ުީ�f�,��:����oE8�ò���d��'�DphDϥH?R�� M��D�Ao"��6������MqElC��g���g�e���.�ՖH̻2D>�P����,�����Uw$���{���T�ۦ�(��]��d�^�k�ܩ�7�gX�6�g|�׷J�Լ�Ѥ����vn��duu��Ifx?����R�	Yw%��W��}/��{�tb�$�i�^���{��KyJ��oG)uр�\㒧����n ���b�޵��iw�!�s)��F�C���(�=/�W�w�b�
� ?<�
���o_���n�h__��O6o���tMB�b-����\�q�� g	ux�� �Z�j\
�g-����T0Y�ߴ<�3̑���{�*5m�b��<).���t)�99JV�Į�T/��j��Y9�g�?����D���߇V����ԧ����ӥՌ"c��Y���yx�� ���!D�Gp`��S�kD����z*��07Z�e��N=k��Ӗt��O���%��P�O���(��,�k��`�)p�`�j����M�&n�X)��^�(�~N2�4�	�B����XR�絃O6=6�ƘDB�z��9B��歿�����T�H7���"�л�IM;��VM��I�\u��T�͒j�Ɇ�Ha��a3��r,c��꼡r)���Im����;���X��H�!!��k1�*�L7 ���C�����&rN9m�WǊ�BZ�{�g� 4`�l��d���:�ႜj�:_S��
8�;L:�-q!S9�8!��Ds�s���&��w����l�{d���	ܨk���d��c>�	�^�
>~�w���T���"~�P�Ԧ���LC�Y�����o�'7[�gx�Ȏ�;y�̆��̲qcF �xML���6���]�}*:���p.���]׀���_T�*r����4h*3�ӯU�ȱ�J.Ũ�� �V��*��<�v��G��N��~�(ꪣ�pS��H�䶆e�ݲ�8ς��h%k���U%��ʖ�h�J��ͩ٫�����<a7�8����+�2:�$;#��E6�|�H�Wo��X��Jo5�c%��my�M��n݅�Ў8H��_7�͞�μG��'C��.�!�2���ހ�J�H���c���e�:��h#����$�/
;΄�x�ey.^��Pq�7�[dl�_V�dҴ����^�XH�2F&���5��f��Ȓ���7�S�oM ����J��.���Y�٠f@�d��45-�q6���zI�
����� ���/��ZNtj(2�*����N�k���a��ٿY�C�p�M[��NZT�]*��d�Hܵ�����[��1t3#��/dM��)~��Z=	�Ī���p�&!�TrD�q�"!Wn�	��<\�H���$�i�r���@�*�4^�gR�ʮ8U���RW��
j��r!�S��O(�:G�_��aӰ���ϙ��F��_��_X������p���R �/U u�ω�F�Z6���v\��>l��2�TΑ*q�d�� �u(2�8���ZX��CZ���)!b)���Ԅ��s�	<J�ou�:xIn�-]�Z-|��);�:�C��o����ReE��f���n	n�%_���l��ֆ�k�u�Ǹ�(���m��zY�ށd`�2:����[�*ڨ�TN�ҟY���8�"1�4��C^��|��F�^�1s7�05
�Z⠂@�U�p��ǈWr��>�3#��o��]�w�a��9���ݓ8��jq������N��ޝ
�Pk7g��+9 e
�4�`�-l����������6��������8���Զ�LO�q�E�e$�Վ��Al�W��Z��=Ę;�h@�Ӥ/TF,d��5��9ȑP���.�%w�^�GyL+	W���ؾ�'����P�����$�_�r�3ˣ��jZ��G�2��:��KN�m��KHU���D�G)7P�i���A<݃%0�ǘ'�"�ME���pu�ES�'l<���o������e�n��z"_���V����'xR�� �y�7��ܰ�S����B8��S�e1 ���ˀ�g�&M��G��uY��!���`Covn!�'��F��MiAU� !���.��o�'>����[4�­h�\l��!�C&��5�[�^�2@���Q��B~���
�-��-���1jұ@H�$)��>������B���GBT':���ehΛ���p����������څT��!:��Q>�F�i6k{� �h�Ra�D��(����Xh6\̓|ʩX��Ҋ��m�nq5��|��Ba�p$&g72F񆋯�0f�73��&���`���	L툧s�C�O��!K��#�lzlUe���>��̡���^�t�ng��0�(�,ͥ�"%��=�z��Ĳ|���-=`�K���3n|`Bnn�����1��-s�o[���hMG^�T���q�'Һ�����P��ܷ#nܧ����Y��u3�[�H\�w��j��sِ�F$�Ο�ԓ�x�R´�yo/ y��~	/#���́_�Ks�(�X��H��d>hC|�)\J6gG���ѷ�b����i
��8M����=���vJ8�Bh�D�����]y	��n��������*g�����w��J�=9~������X>�r�:��ky�߮0=W��6q�0"k����3:T~X���y<�`�$����Yh�%��Iqޝ�վZc� >��^�V�'rƻHy��������v\Ƌ�92r��
�T}�4RN����F��Ư�l���Ň)��q1�'[�%�4ir, @��j�~��'I(��q^F'n�^�*C���SΠ�?����ܽ�[l��k$gQ�i˿6;�� ɶ*72#]���54���^�Ru�pH��kΔ6 4%�uU�*�E/��ގ�3��ѥ��M�a���ߝ+Z����A�!�ԸU�Y:��=e��fW�/�ݴ���lھ^�lsC�7�-]ިt�#Fx�m]+��&��}n���#U�j���7a=��W����|���!^������������/w�CiΝ^��i+�y6Ț�bp���Ǭ���$�x��/�Qm)�?t���J�=^VP�*�/O��
���}(���)n��r��?���e�b��ryb8r���ؾ8���B�-Y�u��#�{h�5�6�nyu	��4�����!81n��JAn�����/��U�݋(�
�^\���~��|t+8s.�ij�2���w-CCK3�����Y5񾼤I��{k�L��z�"�PO{�=�G	���d���>�@F�/73�c�7�6��|�f����]�'�6U�ܬ� b�����J�yo��|�Ӛa?���̒�/�}��55��O;�su�S���Z.��G�>����� ��I�Oν���\.�^Yo��mS�^�����;X��%L��{&bڴx�sd"�V"�QWJᪧnJ�"\��R�3J&�D���]���$R5te1�wZ	� T&w�U4R%"�$4iBVzZ�*?*�z:���:ݷ���o��nH0=_���C����#灞;i<�V���X������Pu��ۺ)��km�P:����D�����؇5Y07C�J�&N�J���σbQ'�:c�ՠS���ݥv+rvf�4�s����8�U�7�H� �����E2Ǉj�י�w}c��Ѣ�+�f�;�7�c�b?
�~� ��i�w�F�[��:����� @@�Uu�
8e�#O�׌N�6���l�՜�.�,` 5�4/�w���4��F��0����G��yi��ʋ�~8>h����\�ү5#'���������[@'�9�c;�*@�0�*� �A >����*v�σ�B��ۙ���6e!�/���.*���+�X�O�8>d8i.3�JFe�x�J������V��Zi��=�YOe�;��0O(��F����W6����nJ���~�G���(M�����?5.���^u�o}$QX4Avq�Ț��c
� �c�V�V݃!�'�I]&Z!V|�݊�k8����y�88���$A�^�5�8m�wL�<_0�>�+D�L�>{����7jX@@r�8oϛ�s��(��/-ٖ��GIkV��@mgka����khK+&�SHE��S��ȯ-�s��w�`���V�	�銦�8C�ay�6ЫBk1l��f����qpDSΰ�}���{]A��{N6�C�9X`�l�2�&i_�n�w�ٛ'�����ڍկ���Ɋ>���|�9�e0dܩH*V�,�@�R��B8-_7���K(I*j��/,|�qi���\#c��~�pxׁq�<"�� &�&�P�t�����!>�X,���n���^��$�ڣ��5�h
�j��8hRԁK@�p,B��r$�B]�Y����ɵ�GXI
�d� f��. ���M*��K���y�G&� ��� U�
��^7��y���
�?�q�2�i��Mxo%+r�WF���y�j���^��#�@��/׌-CF$�Ѡ�k���U����h%� ŽS�ӂI�ҫ�wS�ӝ�8��:��)DMu�ّ�!#�9��8�"��K��FN�]���kz��ǉR��o;�GK com�NUM�HF%	OG-���e`�W��V"�]b2�^���?ո4����'��K�$���+#n=q411�Mr,_5���-z�mi�^��ԟ��e�ŗ��EsG|����SRQ���Иl��n�U�n{mf⌙Ui�+��9!"3�+���m�~��\rw h#�j��[~�7�>��0��&�l�θ3�*�X8j|}O���M�$�ެ�g�E��3a-�dU��p�����s
�!����z��i���	������W���{�=C�@���q�duq��g;c��8k_/�$��eh�A���"��,,���谟�g6�z��*'�`��z�9��$�]J�o��o�����5
L0C]�/���i��g�&8x��t)9eQ{Ys�\w����:쾹���$3�3Ai湜k���k�p=�q<"�;m���	P����:��`肮��dxD���fx�s.8S���
�����ͨ� �q�Gy��±�?A�i�ٴYǉAÖ�k��4���6�o��\WA7m^�ϑ6��U�GW҄�_O�-��J!���Y��`�q*y�����/w=��eoEyp�u�7�R;���ﲪH�(o�7��(5�}��گ�,��hb���4AGW��	!�zb�9͜d�C/�����?���"�'�IC%(�W��s��hEx�~4��>��oe�=t0���X	C���	<����R/��X�Rz\@0���3J�#�/��u�A����,	0���a�Q�-U\�x��/�I�V�XS-b�W����C��.U?w�����;�:�L�2�AQ�@n�H����j�)HW)G�@.��$�.�j e��i8���J"MZ�7.,��y6���#x������߆���ʻ�A��@��=B��sǖ�`ِ�qΞ�:��v��K�����\���7%���X���in´�7��9[�/�SA��g����K{,4}�`p �R�oRD姊�����[��y߆���I���2����=��]��%��w�cK�/��`O��X%��a�B���ϊ�8��e�!7��h�-�'^6lnUy����Y�a�L2Z�	q��w�5;��w��W��jA�$џeİ�F�^Z�c.4�\~	��X=���WWP�
9b�h4G1�mȔ�&(��t��9k�[2��O2�v�6e �8	ɥ���5l5r<�gǘs2_�b-�c���̡ߙ�7�3�v�l����J���<��ap���] +��&L{P���V�]%��H܊�U^1!i��Z	�cv�����?i�='���꤀6�Eh?��Qpg"s5��<�WPq�`����ne��ަ�XE��� h��Uy=>����
a��@�נ�>�'ܵ#�X�Z&�1�̽D d)��y��P0�k�=��Q$�{M�-�u�I��WЎ�����\rB�Ǎ>�8����_-M��ζ�G�����y�4����/�U�F����d\ "IT���fV1NrH"���d#wUGyȍOG��M���4�6��\��?ϋ��\���ذ%����?~8ѻ!F��?�
Hb���3���c����0� ؚ
W�?er��4S\��C�%</X�+�c8Ѿ�������98���|������jˉ;"1��1v��?JD��4	'#���5"��-�okv�� }�vS@����ƻ<� ���	���/�z��G[���ST<R��̷7+�SԻ���sf�������`0�URi�z�d��8z�P���p ��3���lt�&G�U���XQ�^V�ŀy��7���s�LW&8�H��G���b��!<���O����Xj��*��5kbMr}7@w�͹eԺ�Wt9TPw�vn�0�=k�?>Ǘh'����5�7C��=<\a�]y�;:����`fb}��1�b�9�Ň�����U�"�p+f.ZHԷrS��х���r:�ᅺB��N�J��d<b �!�QxY�廸�a� ����WnA���8$�S�4G�y.�����R!<d�;��$ֽM��B�y��Ѵ��e�� ���Z7�ߏM�-$?<˧L��|�um��ڪ��|�hPuK;?������!,���-T��t,��u��/�"Y\�Ю�<�d�d9�6B�?�
@nr��2
5#NΘ�t��fG�O�&���,��X׆���Q-sIWA{��.��O��+L�D>˟��a�e�:�8��n�)h�N\^���vu]�����X�o�euR7=f�P���Mql��A����l�AF��U��x/��QX�U��6Uw&B�QQ�5ɣ[����Q���*�($e(���
��&s����׾�7,��M7�y�6΂�����"�_Sb0�.ѭG�9��	on���Pe�EMS�%��-'XK�m ��_�DC��{ �9S���N�֘l����@�(��d��A�p!��;�W,��f"ڴ�:�a�M.<� �D��˹
��&<�8;Y&�v�R6��Ui7V����y,=\�R\] ��f�z�m<��j�����p��IR�|:���:�\���-�U���Y4߹ ����9�����%�{�<�ڗ��]X������,G7/�a��݆ᖠ�b�;�wҗ��dO�ч17�{J�ex��Q�s��+�-ۧ�۫�,��C�m�_v�Kӕ�9��T�HS@`��wr���<�֘��@bU(�?�k�"<k<�]n���k�5-%����>M�[�3��h�x%K$���������?�H���s����Ұ�V�Vە"w��p�	�K@LRzϰ���S����}�C���_Z��	�s���#�wk��k��`��؆T�up�F���(�Ӕ6��H�M'�1�-զAz�Ք��)(��o�ZDp�<[��u����.�1�CUQ+;�Vq�b/�Gj����]��4dV�v�CA��)U)���tGҀ�C�gf��cw���u�2"I�4��hQ�FM����x�CҼv�|>�  ���Hq��t��՞wſ�ߠ�8�] \6&��dg��b�m�aQ�rb5�J�Zhԏq��mʒ��g¾����TK�d%�jR���SV8.}�����l$�D-}�������(���1tpC�J�/q��ҫ��<!6��wg˘���{[;'{޽�hxb�4g��z�d�o�[��_�̙��6M��ݵ+�<���z��Na���N�{@LW��_'f�(rn�0��OR��-�Nn����p�:|L�ج�\<
�x[8L��u0_T�RP���Ar����#��m���^N(-_��[�&��l͈翙�6�W�N�����1� ښ�����.�BK>�X��+���RX�b��
���X�p���yʃ!3����Puin�,��G笈x�UJ$j%�Z�(ۦD$@�b�23h��E�h��\��� =�O���|�Y���#�F�{�t�4N����@� �߄m�;��\ ���vB�h����䶩Lv��jW>/�pt���s�A�T�s��\j۵W�!I<�J���h�re�OsV� {w=��?T��'�-��9x]$.��3LsHM��O�%�hL�Τ�$\�Q7b��� B�nS3z�-��!R����!�s.����'������c����sedQ��/%��1k s��`3/� �=yǞ���i��Y�oJ�Z�B�����Ă�������d'�r�J1gk�LC[=�ࡴ�Z�s�p#;�g/�Aʰ_k�Q{	��>�[�Th�0�[�r�W�؛�k������L��(�<�l(���o�g X�U�Xg�xSCv�M,>-�;ݕ��V��m��D�ée��aT���zJ�Eaŉ#p��������杬-o������2��>bM�����T�����)Ȅ�RQoD��f�t8��ƍ�Kx*�k�C]W��n|��� <�a� I6	%�P]0e�:�%X�M�gsTd/��0�x����B� �����K�n%A �o-�V�$F��.(�k�\_w�1�=��d����,x�(z���7�dn�%U9�R�	�S���+v�9�}S!��?�i1o��0�:��qA㑸#�I�r���7Uk�<��3)x�Y������X	DP�0�&��E]��"��}��6_�A\���{ �n��/F_ܴ%�RT� i�j�]�$_���%�t��HLK4+���G
)$ �1�:�AK�Ϊ���3���Bțjr(�zPg���eP.c ��dla��9C.sGݍ� Rlɓo�g����xH���^�
�& `ܷehC f�J(���z�� kXL�8���d�� ��*������}��ْ�F�)�"�e��HK誦!�X��4��[h�9.���.R��K&l	�5i�����5ݫ�ӥ�8_�k�8�1?��峌6�]{V���C*�ԓ�W+�OY�B�l�]&}���ၻV82� �����C��{ϓ������Omq��ɠ�����5�>xΫ�V	��d�����tw�Î�U��5��ǾXU�>��D�����o[VB8D�/x�fqe[����d%2������V����"�n�04d�_*A��J�FN�Y���шr7VAL�1%`��w%��9��V�,8�Ս���ݲ�� 4�*bD���a��^��c��pֿ���FV�K0�>&�5�f���)�M0�H)��9D>�<x��ϮܨK���:P����f��W�2^8�j4]G9"gn��Δi��nJ�0�Dݭ��J�����s]��$76q3P�^�˚���@l�&�_ҀM���a�#�9+���U�8l�)��zĥ������v j�-������tY ��T�V����D�B�/���%��a���RT��.�g���� w�A�G�:Czߍ��`d��d����Z�`S��IKfU�^hإ<�5xL/>��� 
���8|�՟���a��m���ˑ�Ş� q߾Y[Rmk̘;?��d�M�|���"$I�cq|%Ҕ��Sz{+'�?�j?v��\N$j�^���(�H/_�\%�x�x���Oi��s��\_��H�rd�½P��x�Т4�b�CPg��*M򅵆�g[&ug$������6�'�Ib��S�+�4_������C�~�L��l���&�������E!��!~e��h�,ƕ�z�X��Ҝ�1l�~��{Q���T�/�Z0��mG �.Kʍ������ۿދ@*�����t���-�����
�Ѽ^�]DiQkKsAY`��B��u�j	���ʆ����w"1y0�mk��.lh����jR�t�s�lGL]�y!|����¤g=�WW����eK8�/�������HL&��Z(G�x�n�%�V�̭N�l||� =(@�����a��|��S�E����_�e�%|m,���y�|<U�O�V
�5���"�С^�蹕�R�]�n,,	� �TA��Yz�(��Ah�[ɓi+
���I�;�֯7��v׍�o��~ G�}�2sl{?�C ����L��|�G*1����7⫄�Q��Tt�T�� �Ä�?��:���14w|��O�n��A�x@@����y8K�@�-������l���۫�*ݠ�i9s5ТI�9�z�B�繀���d��E����6�OPB�+S\!Q���A���]���8����b<��j@g��>���5% �.@*���T���d׏�F������.�Τ8A�����ا�aS��Dw��{��2�X�E!F�[A
/�~�8�Xj�c��F�
ע353{�!%�YS ��oi>ݎ�Z@��N	��;�������'d��IB�떏�����`ن���W�׾C�+'��(}�#Q��"��\9}6�;g�Il��s�#ַjG �@����Y�3P�cӡ��L/��W��+���������Ej��T��3��5f���fs�1�ڷYVTvJ�0z��` �B�4�ɋ��3s�j+��D)�:.T�Ѻ������o��33�N�Kk�G@�hV��s¹q�O�E+@G��2�-���߶U���!S;I�EI���WӦܬR��^���w6�;q�i$F��"3���N�j���ගu�XF�x�&�G���_Ӑ��!]����+�}C�v;w���e_y��;B�Fk���ڽݮ̑�n��J6�	_$�ue,:c��1u�yϧ�k�bo�И2=T�>���Z�c�����߆�8�2�qPPt�����M��<��j5�����.W�R!ns�c����l����j�4�
k�6���5ٻXv�db��|1�G��<]߄�=o[4t�b�9�Q��p)�CÃ�C��UR��x)�|H�sD*�$m��8	�JP��E��cT�����~��=�b���D�4�k��ᴻ�19/2w����^2�p]�2�'2���|�ak��.�$ꍁ&m��:Q�1�4���L<��&g�:9�@�bS՘��0�fL���>Q�5�ڭ�.��A`�dqe�J0�ࡼ\��Nw���SX�FㅬV�@��d�+o��7~_g�@l)TAy���9�$�HG8�u��g�<���m�z��a�
ŤC��t9$��m3�-�sXְ�$�n��q3���d;1u�z��:�\�����j�o��kJ2���t����S(ɑ��}��q��o��$�g[��~�z#j�Nrj*/�KhT����Đف4��z�����B@�>�-����B���NN> �|�'ym����L\$9����@yu���j��X"#�}��{D�V[c�L�-R�}�"���"��� _6Ɯ�R�F�jIF��FN�(�d�=���V���-UЦx:G=��ʊ����A�����{�a�$�}�1��"kc��yǺi;̆ڙ��c��ѽA�ȣ�Lb��O���A��۸Imn��%����x��]4i�
�Obg�ȓ_�e�_M+����Gև���o�cT.
�Ë�t�a~���v�=l��ُ��S�����pw��M$Q
}�@9'~lHt~���0�^	�2��A��!����F͑͵ٍJ������N+{�PU�ݐ*�aeOL�s	C(�_�I���4@�d�/��J��y�9o����B�5Sz[L$�#�w���~js�9�U#��J�V��f�sX�|��&Zq;CX>�t�t��G���>�޷��+`_�y�N��Akw�;F~�]O���㽚�Rϫ�?�����N�j{��|��R˜-�G�Ɔ~f!���M����A���]eB��'Y���;ا�L� ���s/�
C<��	}]E@�5n��h2�����j����;�ѣ�҉f�L��U�^7���z�P�J +�x�X f��!|�&<4l�J#�x0�=թ����:� Xd>�KB����Ukl9��m�"0^]��A�rJ)K�e�*�������i�q�oa�(d�:���L*�M"�>4�adU��i����DQ�]qH'*S;�d�8�ۀԢ����ʅ�3r�c���E"T�����K�w3�E9��~���&3�LC���O�����o��N���{؍΁B�w ��T�y">��$~Q�g�lzBV�?�1}����������~����!X�r474�M��֙�c%�J�T��[hI�4��K�����J��Ι{����%��_�:�L3\B업J�O)��b
�	�a�&fNP}�';��pg
�ob[p�c�S��'���	XR���ձ��.T{�f�%�{ts��u(�hv�{3@��pQ���|����B�5���5wD�E�U��S�m�l8��|�m1ր�H�
ҤE�PKϸ�A�n��y��c���\z��ֵ[3Z&RS�2��Й��Ei���Yr�>l�,�n��L�;� �5$�I�b��~mV��S���["�&�.�>7j1?�C��b����9�\�v�C���$�v=�[`��L�0	���M���� z�g<)o#7�H����u�D�	L���}3���*3��`>u��e����/[�������ȘT���w����&)!�sز"c����>���VH�E
O�:�ao4vB�lQ�j�m���0�>6p��p����}�T?F \Eqȁ�h\�H��{ݻ҉�����+���Su }mw"uR���w�+�,�	�<�.==����,ΰ;C�����9
����O>���� 
�&3�������ӂ�猇���.�Q㝾�O]��C�d ����R�oo�̀�y~&���ӊ�OFM^]St�9��&���m��n�>�F�����v�Y��֌�0��Y�oT��M ROE�`5��4���}͒��)_>~ݼ2��\����2v.����)��|�M�С�����ed$��~���~���AXrg1�?̔��i���d'�~��]��� 8������/c�y� ��(ݼ�ĵ�R᫋|Ѡ�vP�����ȞhLVY�!Ԓ�a/�A*�{s��]P�BG�J֙��p��a+�Aca��B��h�O���P�sl�	���"J��ۀ�9O+y�d��
%�v>6"�� Ȼ��1�"���_%��S�ֆ�:}|��=u$�����{��j���%Z�k5���t����[hw����\m�R�jr(|Jˇ�1�tܿx�e�u�vKz�վ����ߥx�(�Ug�3��QO��X}������h{U���	�MCj"h;�X�qP<e�~L�@<p�og�n�F�T��
9����;�M��ʆT�t9�-����x�=81�i0q�z�$��h���~������:���<ڔXdц�&��2��<�j��՟(��F��z���I�3?���a%��h��ס~���8����-$���_B$��E�I�/I(흣Qǯ誓�h<��a���"��:���׸@y�Q�06`t��^�<�S�uh�9!�6�}���d=z�.g�z���e��3!y{M/��_:Z�Z8܍��g�Z~�JX��L�`v)U?�Z� Y)��#6IϟM�3?�E|*��%������pUSf�ّh��8B�����<%Txr��^�,�G�)*v�C&;O�ޖg{.y�� �7p�o��f�!�7fp�cE�!jn�0������G�j����K�g��}��X/Ο*�N�Tg¢ ��'f[��[�g��ۿu�c��D�"N9��~[�a��>�̀�b<	]��H�Ι��D�dcߤ�&r&6�#F�La2ްNy����z�������=ҍKM��
X�J�'(o�Zd�}�/�C����;yzB|fHQܠ�f8�&X�|�����g2M�χOfd�����:�(`bR��Wl˨���B�0�$X����%�cIG6[��s�a�%g�~��`��|*���z�~��$�8�����:�?N�aM?�J�%�����a���3N���)���5�(XMpыv!��X�Eg�v�-E�@9ɰL��<e#`Pc�)q�dݻ� �"�������j�T�S<��H��(��� 	�9g&p.� �S��<c���ݸ����. ��@���_&G�q����h�*O���[�ϖ��T�r[Æ��_x���t�3�>#��t{�*�U�'͸	`_H�C�	��x��j9�IO.����i��i�Ї>F��9��/Mv�1i+h���\P��t���hD&��Uˋia���q����@ r;}#nS�5�93�eN�]�&sR@L�U�o��j�@D���L���C��J�l�'A��g.��U�#�N���9���i���|aAX���FjnY8�g=]~ECE\/B���R�V6�ւj���OǏUkE��_p?�g\C��8?�]Ȕ�;�{hu2��N *C�uG�B&k.�����i+�բz�b�z΀�Cx�['��`�HT�2���1����"o(�o�h�m_��(0�!涢K��9�C塉ڕ�Ճ@h��ߥt5X̀�`S�����?X�GFN|�6�׍� M�#��칸��5v`\��~�����z7ͬ�M���"7x�����;��ĐV�*�qgVI쵼{���K��^
"��V�Ań��R1#X/8�y�|�O��x��5P�c�գ15���d�
���&���%�y��Q����A�ͼ�up̕��^����̚���A��T*B`���p>���!)���r�Aɝ�����<���pR�Tŧ ǳ���'�񁀏HΦ���vX�iY�/N%��s?��ţ�����C�N�5ė��r_;���5��I��=(+�	�n��{�{q�	{�>,�=����� ���������*�����h�p�T�g����`�{�7A�r̷v��sKf��G���ҥ����}��o����K��?�#N؎<��á�i�X�����8������F�R-�t[hJ4 U��b�<'&�Dќ�b�o��|�h�>�y��c�2R��̽�� ##�Y��?�QSS����/fVA� |l�V �Bg�^hٜ��潩��������j���s�jںA����B�䳡x��lHK�F�y�E}�k�G�F!�=}�;$���v���5�L��+|����%1Om��ρԣ��S:b��ߗ�1���;I;TϏ;��h�3a��w�໸���4��^�T�PT�{� ��>5
,��W��WB鵙��Pǅ.��
�_�&4��?��x�`�PU�
Q��ۜ>�}y ���(9Sm�d�Yx�����V��Q����i��J�� ^#c/锘���\�-�[Q��D�� ��?hy+�������~�Ue�Lǂ�|#�7t�W��,ڑF|*���\�Q���N���oS��q�>ň���2��ZZ���?����Ƿ/&rz�#� r38�R��|�#�P�y{���I���yiDD-��Z7Q����8
d/���&)�M	LQ�/� ���g��d�[1Ҽs?���0��R����!�-�T?�^#S��V?�-���5�V��Ro���n�����h��l�>,&	)��B����[�3[o�������_����O'4%{�m
k¶?;�*	�`��*!�b!%H�F_���Yޖ/Rz�fmN[�F��z��[�ۗ��lf�[���qe�b��IyE���t��f��WB�o���}V&�A�1>���-4>PeW���wK簕�p�)�WX3�{�
�=@�Z�cy+N�����H3>����24d��o���_�Jn���V�'��U�52��m�\��"�Q}�J�4�@`��^�w�/7�NRoAԨO�5e�΢D���������y�\�F���T�_Sp�5~�<4�<�o:���:��k$�� O���52��ӊ�t�F{;�3�h��%o�mrYt��h,�k1��`�yzP@�}|0���$���h��<�1 �Ie�WѢ�+��1�c��O����8zU$ ��=�8o�u&Wp�=�1Nj}�2���|���g{��%�ʦ?j��6X���c����+��Rz��6�*�dڌ�:lI�>��m!������!�XT�\=�F�X��؝.�/%(�w.M��jcu*2I>�1������VB�~/XFJ�C��;���HvQ���h��)��H���7ņ��{��N�
� ���_�X����a6l�j.�W�� �[CA�>��<zg������*It=羏q�;�
���<�n�����,��f�Q���g����z��K{& _65��=[\%��AK�<�N�~���$�W�B��9~c�5b}��^��H��J�k��4t^���ǖW�����F�	mU[�
b�F��y���[�Y���u-�
IRz}\�T�y��1�nn¾�z��+ ��{e�@QV����.)}�ŉ�ؐ�r�Tt�x�g��y�~�$g��	��z"N�RB�hj������K�2[�Q�s~>��DP�k-���<��V�N��Ʈc2`�Iq����W��@h��'�LU6��˒׭(���Z�:�$�}��0��9�Vs�Sa,;���<؎ I�� �`a�G�Ʈ�?{�(_��ѣԄ�l��_/D鬌�yRj�Рw�jQ]o���~�� ���'^3D��g}�bcLv���׋����R���)b��ޤ�Tת�D��@u�*[�g5�ލfR�&#�(C�c��`��v�;wN�����pĒ��w�b^`�d�9�� Gk^�I�jvf��/=[[ �bm�������Ѡ%sX����އW
w�ϖ] ����$jt�<��ۀ�!YZD���!�M>��0tA�xw��K�SZ|�}���)�L{6 j����v.F,46��q8`[)
���nY�+����x:Y�L)AJ������������$~��	xC$n��BE�9/
���*��Q�S�/��/ �@I��r���3�YJ��&`���: ��3�4�=��
u��&XVNPޥ�|,�!���Nf�s����uͣ"�d����FQ�m���S?@�����j��a�H��m����E_.OHH��_o�H�yy9Jd�8����z-���kH|���	��no��i���1_C���,�Ǵh��~w�i�%�����d�q8hd������O�u�0����>k�a�T]��
��|�ҙԼ�/��?�[#�?��H:Yև�)cٹ����W�` C��Gu��m]�.~'���
8GgtО9�.=�������m���V���l������2��b�<�^��J-\�.2�讏��D.`+[ձ7�w��L�8�4~�貒�S��J�^SȪ#^�|�rl5�D�8�.�ޑ��Q<Q�>���|��	I���5�-�9���H(�NN��>��&PU�?r 2��k�|�a$8W��=��$
��~�	3�ُ)r�V��a�m�D�=y%�W鱩���.���bH&��+��*�liz��4źx��8|��
�������U��(�����/��HM���!惫�1�Ni=���넱l���K�0'T�9�+(��;<�qaE�p����LX��Y�Q�����1Q6��|�i(����x��4N"\�QtW��ю��� ѰLD��G�e
)�����D��L�x�]�~퇌�*?�F�;S}����=�>b�����R��w��6����D��""z1?�fU�-x����i�����.aJ���9؝3:.��L�
g��g��s%r����	U�ZW~�G��:����3]i�6R&CJ	�s�J~�������X?G[�jU������6|�O�×��xG��7h����,��Er`#'�`��:�&e�q'x٩9q���NɆ'�3�3J�橤TkUM�
z�â�<� j/Ě���@�{H�hG�%��0;~����a��i�%E>ϋ��;�����F��U�/@�X��K�yG<���I�Q�Yl��H��&�&4Z�0X�2����`f��k~zo�E����kqkI�u��M��L��EHo�r�D�xJ����FnxR��2�nF�����z�2,��W�������T��z��j�GP&'W{~��~��br�*MQ�Y�Fj�B���{��w�j�ʶz�p|l
5��}jϕĻ��DٖG\��	�G7T����'+]_$�'��s+�`�<*�a�poG�x�IT��įn��::R��D�w�-�Y������]������;
�����M��
L\8J�卤k\�*�p�-�����\�o�eE�6����g�u��f�-��<L�l�_����Q��n&���.�_ϡ��6�5;=ӓ��:;ɾ�����L��oP%�.I��vV�*j�%!tV]<�����АKK�K��m�1��I�t+���nr��
Ao�7�U���h����x�Dw�cgG�m���� p��
�|��y�r�?�Cj2���eE���At�'�$<^1�#N(��&���0^f�%N9�j�<��u�'/��i{jy����0��w�G�a��T|7�O�I�5!p�zʨ:sn�������)pL��5��Oʪ�xIY!0�oac��aE�H}��q�����n�4=�>_M�ko�3��E���?�'s��_��Jg�}�����h���o��%e6u$�_Z5~b��y�Oȱ���1äS99�ʑѤ���?�<���~�2����7P��ʽ�W��	*��'I+`�;t]�!� 2�O�(�v��ے̫0�:u��{���5W��:d�23�Vz����v��ck�%�;�.�����Ӂt�P�Q)k��g;n�=-��;���p���kH�X������X�|ܽ ���]@7k�.��ؼVoh_Ji�Ø���q<�rs�v�Kb��,����M�?� r�Cr��i�<F9K�]�� 1ć)�ꅄui�3�#��B�O%�Ӛ���V|/��r��y�(�opT�M�h�H��<~o���w���`�O�$�T(4�,�Lf�B��(]js��Ң^����m��}#���~k���@�Ҭץ�-���H�8ˮw��Q$:˳�!y���-��P��󻘃=�N�\S�w���D;�S���q⳽ �GP�N}b&I%�Y�� V�)O���w��n�LI�倯.09a�t�7\%�s�3j��W/v,@T3�>M�E["Wn���T��B��-��U>��~ү���O��_��p���#��������]0D��rd����*��Z<o�T�<����vL����Y�AؐU@T`�ܺ5��D�G�Q[.���^7jƻ�[_�w����&���=����-�͆�����`��9j(3�-*�ޔ�P�b��¶����f�d�vw�ӆ����������Y�f�\�A�uR�Xs,j+4��N�K����8��P��at�^�����ê�=�.�ٽь	�B��	��x��`��^Tޯq�:%#v(�L�[:�g��o��hX
���Ģ+�ikg/�PZЙ45���L��<����X������Flʂ#��p1J/��  �@��
F���k2g(�f�O�Z�����M�1�o���Ŀ�LS|����ZG<��07|��i8ǵ_:ז�/.*݉�?�c��4��u�4U�i�gn�sHǈE��\��IH_	V��P�_�Ĉ��\b4�W�H�}~��3>^��I#%h�S�=Q�"اw��������"�����J��ojֹ�uR|f�b��9���T_���H��-���y٘	"�o�&��TG�4���r����	�<ɛH���ge�B��n�wi\v��4;x��p̙Z-�����F��ѿ�s-�#B��TO;aE�xA���	�y�jXC_%���� E�l�3@t��?cj�`In&x�k�Wš��a�Q��c=��@��d���΁vw��g�b��Mط�Nv����ƶ�󉈪;L���s��1}B	����q��#����1��u?|���3�fj��܁?�b��	=��r�O�B�ӘXo�:�����C�n��&UUdp�
�<�w��R��%!�qX���
w�Ь_Vo�/]Ӎz�;��s�?��g6&�<0�{?�ydO�M(���ϑ|�G���Y��W��[A��mVFA܃��<`̺�1V=���|׺�a݀6��{�T��t�dZ:hH8���z:������%���;~~ٱE��??�`��'ǡ��׿Q�����$�����[��{ɰ�7gCZ�&2���d
�I��]�@�Z�ݏP��r"�`W�>&������:_>}::�Sb;ж'�:��e���{M����;GX{��6����삳�At�f�	��[��e-jJ}�h��e$��K�v��外�ѯk��?u@ژy���Q�5�ꢊ�h��2`�5]v��bĞ�*=��Ѕ���X��v��\��������4��+S��g���u� ܋4���k�]�~����Ƨ�v�x1�����+�~j���ӕ�� p��T�,�� ���d��u�!i���*n3���E��R� J��0�`Z��p:Ӌ`ќN-�SҎ�Y gq#���sy:�j�ٔ�C�V��Y)i�B���J��0Uد�V5��{?��Y�i�vo�^ӳ�f�Ћ�Q/G�f~��R��l����X���L���	����y���/ml~8y[������%;��|�]����[���g�O6c���)px��͕o�q˿�̖ d���C�"ү�I~�ʣ?E� �E��I�&�����������C�+���5}xD.Y+j:�Ycj�L�O
v�YՍܸ"L{��w/Z*ʝ�\d�<i�=��>O�pCy �ݏ�k�ew��pV�D��3�tl$+޶�#w�fΈs~ɞ��+�6 ��^J�Bk�h�������ʚ)vD�����o����dW���l�A���#]��/�z��t�p��`��G9ݗ��ɫ��><��&h�d^�Ku!��݉^����ra���9�i�[��'"�_����݅����ϡ�7M]�P����Q>\V���E��>a+��d�� ���j|i� �8�?��Fj��IKF}�Yc`��ݔҩF��l(Yv�N؇�緥���(�3k���W�|J�(����wG�r�_�Z�`\�h);���P���6�j��(��d⦓�&f/����?���݇?���dp،��WA��T���D���,t�a�Y$!i'0��ϊ�05:�0��\�� �>�mܸ!��=����?��7� H�lz@�iR��|!�(EʀCZ�P�Ҭ���3��n���Q��yn���?��ߜ��l1=�$�E�j=,�0zy(��.!�V���x0��9j
��w�X�9���y�z�%�v����?R/Ku��Y��0�j�M$�]�]'�zy�����2�Rznt>:R�/1�1w۪4]���(�Nq�ߑ�uX���b��إ���:h��q&D�on�!��� �"T[��p<�;[y���U�>W�P�r�}���ˏ�L,�.2ޥ���V���}��{?���k�MH�d���bH����M�x7BA�SK����8�a�۹���]~��Y�X̊�b�l:cKЬ<@��E"%�H�Y����Нd#��1gEr
�w

��$��E�2
i�Z�ӑtU��׾�4Z}�J|�I���\��I�:�M�$������fX����ib^َ�br�J+wF��i�/'SX��}�u��%9�Z�b�-��|=ۚ������JC
����"�M�Y	Lߩ�P�y��m���BQ��Z���.�ˠն;F��rb��Q�,VE�`�f�*��L��zȝ"߫���w;�I�����g���H7�l�w���$�'�	��c�Gm#�YQ'Z�s�Z���
�s9��	��F. "۽�@�l���ȱˊ��P��u3���+*lUA��?��!��6,by�[@4v�v�ˆzo�'Jql�+�U+�rCK�i�a���a���7E�&�]Hs�ÆS6#.�̓;�����`d?cOHG�?7T� $G�5��N8woB%��qB�p��hL�!������������Y씁�4c�0�1);��:���?/����J����uO���u��2�1G��$��h�u,�R ؁{3��''�Q�������zIt��LK�KUmLQ��U�%J
F)H���L
S#�+�2���W���۾-X��%	�=wj1��.��<ZG��%{�2%��s?����:OB��I�z�LNt�C�NZ9�M���)b��=���X�.x���Z:�:�A�]��8���*[W�u��Jc�]~F���h��<jS����QT^�>�K��J �Α�O���_�S�ll�F�(����%�O�Q��b/� �	б�R�oY]Q��t--�f|]&��%(����T�R��;!�M~P���/7���
;ٷ�:�5���))�����T���C��:�~�=�!�BVY���wZ�Ȍ;7��qiR��q��(���^f�V��o���QW�����CΎ(1����xJ�rI�����ZanF7|��b#(�_C�d9 �|����v��xM�`��������KA0��s8���83��y#T/&`y
�Z�P��E�{k��y̱�b��(?�i�ۗ��0��~�+��zM �T�`� K���p"��s����'�/�d��C�^8���k#�M�Ć��V-A�.1�cC�Q�W3���/b�)�FO_��R1[��-�T�)&w��qҽ��+x*mG�p��������`���ŀ54�'��Emt✶��,��1
��1fw�Y7ٟ����)Z.v�wږy�䮐�?]� 6�ZTC��J��c��H!z�)��-i���}զ��u�$"��✁?�cɥٛ2@Ya�+ ��+k�&�tؐ"K�Z�6M8�l�FX��������o���.oT�1���.:�l	X�ك��$�AU�ײ*1p��f���d�d,8��'f����2("0А /Р���l��,���9A(w����@��d�_k�%���U��CĐ-A�KK_�̴b��=_�V?�^�-C�c��HE�L�5�&$��|CK/{=|e5#�:����`;YRӒu���_ �9�k�R2"�j$�˪�*�t'U��
���b8
	������9|q,eYzu��۸Da��Nʝ���S1����p'*�b�ͫ��}jqd����̜  �I�yW�a�6؝�mc3"�������H�vH��}w�p;��qʯI7!���dh\��ocM�ؐ�ng�f��Ͼ�0��M�IQ�\*A�@eXb���Z{ؘ�i|}Q(��3��k5͝� (�ͮ0�6������)ar��k�D�b`�N� |��ki�#�7��� �����e�c�İ6:�8�>���_��/��J ~��[,��B�C�V��
`\ ��ע�;^�>�����Q���߭�`�4�����fK�GG��Ç^����U�nUB|�oNg�}�o�-G��U��ʎ|FJ�;�1�N-��=��\��>Ylfg��o�Ok���婸����
i�YdןJ�'�Υ�f&�����Wls�P�rًS"�z�Z�G_�o�����%�}7%]��H�R�%��*P���4�=G��ǵ�OI���f+�x�Y���X�=1�)���z�WU��
�n:��7-��PO ��R�q��D�X��'��Y�΃a�FI��]�/����(�_޵s���)�(�t���)a`����f���.��?"hck��a"���҇<U��hX!ə�MQ�lf�eV0^���$���A���} ���^��@n5���%��x W�.���?���`�^e���uU		��da�,�ǃ�؅����A�:�OՉWj��x�Q��o��X"w�ͮ�R�Td2u[���6_�Q￢��T?���=��j�v�\l~Tf�����q9��2w���}ʪ�7;Y{�\�"�@�xc�I�c0ѝL���@�BU�m_�Ju�\̟W�)1��)MlA�!���!�J@�n�2�I�6�д�t��&U�TƠ������	�o�d6�j  ��i��6��}%m��sW���xpz���W��+Ƿ�z����Y���nx(Q�^l_�
A���O�����_�p���"��z�UR-�Aa��D���3��@Ec�R�`p7X6��ji����I���<��4�ğ��}xHO"�
p�j�n8%�O�ܝ�Lj��-'�3�q��Ai�G����p���Yʴ!�W�����7Iz�����?�N~����f��bΞfQ#���a�\1$�ݽ��	t��"¬6�� ���J��u5=����vP7�hp2�q9H'5IR�RN�ke����nwD��B0�G�l͙7��D�8 �n©;�^�-�I��s�g�/Z�J����K���wm�W��K��~��$�Ͳ�;�H��z�PM�&� }]�u��&f����o�
%��C[V���ش��n��쾜������
ɿ�C(&��m
Li�� �&#!Ie���"Y���Ux
���>�qz�r[w¨��BO<�)^��z�X�;�s)�"/B$��y���(b���Z����<ɑ���'y�����/0wx\E>�Z���a���[�OO��Me(,��P���у6}H[�r$��,q�m�"Q�u�	�s򜴮G�|z��ͬT>��ʐ\i#��]z+^���Jɝ�%-�^��P�EHi�6t. 0��j�`SV��һav|*kg`�H�w�!3���Ъ�t���|F�_�8���vC;��ɻ��������(��X~?����4|�sO?oT�iP2��U�{���P�Z�{3���}��N���H��7M�b1dHQ�����3x���x\��M��G8�0G���Δu	��7	�_���h��LAHL"�����-t�x?A�n�6�?Y<�L����(A���!���x�$3�:�������I�y�3���p,�,�힘3��x�EB��r��? T�,5���f�(����ܧE'��4��s&V)�x='�-r���`pq&/��Ҟ�!`�(O��b3d�l�iJ����\�|�V��s�/�2��TMW~$2�x��������"�+�`�����Tws��O�:�蜷��٠���XM1��G��r����y�h�e�^�Y�<l�?��}�Z��F��}I�W����RP.@GJt�q���<M�H��1h��E>�\����`�q�j_d��V�/|:VDL��υz��)qx�K�_2$�?1��ɍ� ������j0����+���dbS8��8�[_5DG�RCưU�6�5�~Ŗlg���O�[�cꂊ�4��Yc����z���d-v|��V�s��qQ?�;�]�Ҩ�Mu���������	�9����q�o�%>Ef���0A� M�y�О�j��"�V�a!¾ʥu&��38��{3�w���2�y�L�_��G�)r
�u���'4;u���k\�'���ΓϩV�7�*@�a��*���']-�W8x��[�kzw0���=�O�وKS���pJ1�)I�ͭ�&���F.�4�T�j��L��qL�7y�a�CϦ5;1�@o=!�3�x�#��NJ��CH�m��FKX�@A��[�h���ӆ�����R|�w�2=Y�Yru�Lu�A�,.�Ip���V0U�(4Xx4.��ʈ��G���.���x�����>�9�d�g��������[
,�8���#�y���b�z�id���ũ/lm���shN��� ��tX��@UC��L����$r
�"F���A+0�fg��������1����-k�L��"ߐ+x7�:�HkKò֚�0��I�,�l��#8F������+E/P�D�ӻ+�E��"�]�����I�F��l�WM'"9ݘ8��c8�QB�S�[��8��ly��rL���:�m�6{i���
d"g����2�������+{��m �|?G@Dd g���O�~����t]ŦL�w㙱0xR7�ǯ��ϠfE_��7U9&���l�Sr���RŴ���w���l�
�,�Fh�;�_n�,�;��1|�y\
���Wi�tŉ����7N&nO�d�5Ż��C�tu��Wj��l��,"����p��V���<�����U
Ŗ����Y�Ӧ�IJ�#����*�`�0��	��dЭ�� T5�8����ҽ��K�����T�I� ��wm��p��ԙ�Fk�\@����Y��B�����C~ĹL����O����_N���\�O�F�N�HT}�/�Hƫ�sؙ�+	���ya�����S�?��yo�,�w4�0��#ʤ ��*R����Ǹf*��:"{�-&ll[G��@���&�oT�^����NQ�x����r���%�n�qX]��{5��`��EU0%]�$	z�sZd7V8�}f�Q��9b�f�v`S��E�M�R���p(���f��� ��_����T<���7��9�/٭���
 ץ�e�T��?*�NO�����a�
"ba�4e������ӝBZҾ\i��\�a�D��[C�)
�s�; �����.T[-�ZP��=��g.実��&��o�`���1ihP�����EV�?�:��j�z�CPx1��jj�����I�!>��3̶J5ޢ e�*��qP�q�:[sD�<���t/���Ԣ.y�M�y;9BU���K��OkBc��XWB�x<!��-=��+�\�p�I�w"���"�qeEL�N۹�b�Sw�$xR2��Q�̡��zQ0K���/Q��fi�a��!FC:�2�%�K%=9��LP�u%��K���*�nE�Y#sen��M3�r��������W�M���*�@ZL�k�o�y��������GU0�H�]���/�o������\��e���f�ה�ĝk�2Th���᭣*�H��3�'�� >�"�6��"����oe`��\x�� qrZܟ���0��PU�d��]����L���E��n�BS�}��b$���ѷ��V�%d�2`�e��<��ǃ%n�;�[%_�#���Z\��Z�@�������2�����Cc�nY�DRۍm���W�'B�:a{�� ����2^�G}:��6�$r)�z���[E��|�A�W�<*q�۠]Q ��R:G���m� #g��E!N
��k����yy��JE�A�����^�>�"Ը
L���.V�{*tW��#2�ͅx��ې��P��o�j%AH'm$Pq	ğ�]�Ĺ( w��*�-V�p�Y�}�3�¤�}������1��Q�X<3F !5��l�p�_��<?j\3��I� ��κ�:�s� v�/ᝌ�xXË�>�%4*YY��'�o�����M��Ԗ�f�j<����O��.����^��Ǉ���e܈����Wj��'����iQ�$�{����R%�\aCS ��l���w�%�n������;8>{�1>��D���V���YU�}�}���� g'p�f?\Oׄ��D����m��t+CA�³Pö�t��@*w!��0*��<�?o>0͖\�m(���͂�a�-cM&�S+V%��J�@J��1ҩ�%G������@.��� �4J���*��P5�2�7@B:�. �w��Ƽ&����Lԉ�MD��	5⩿�%��|.?U<��x�5Z�ҋ��\Dv3�XާF�Ű�9?l*߄�<{�����TH��(�^y8a<�j~y+�ᩏ1����D�:_�VK�(��&�̐�tP`b��YH�.�M�~H�8�A�x�K/��I��\%G�2�8�+̺��T���m;*����������%��z��N�%����t����Zf[�eIY�3�n���L�&6��p�pX���x�Y(n�Y*J=io^m���Z��$g��-�ȵ�Ŗ]�&�5�3	8@�-�|�'���f��nsA��k�:c��,���n���*v�K���±���FQ�i�ps���~�`�.�N�������8��85J�ii�s ���;I�7�K�8W7��	ś��#��f�6��UnC�/���K�~��7h������z�Aj��L8�V*�±�Gڛ�T�A���<:$n{6#��5��~D�O�`�����'Sq�vjV9��Hz$� -�T���FW��"p��X묖��v���=�7�ô �L��s��DՐJ�_%g��=�)��L�!1��kw,rE
`����O܉�c�,87�Uɉ̐�T?���[9l������H��֕ie���9�����C;�E�c&+B��&+��w_��d��V���_(WI+Z=cL�PI��c�
����=HB�Z=`�V��7Ha��H�B��Jڱ�ւ�4��O��D�;O�����h�4��om|���.C�Rq=�R��P��Z?��R�2D�@*�8��:�MPxkfOA��[(Z~1~�1P0���C59�_oԝG��z2��nO��ν��T��>d�ۄ<l�W��-]���/�E��	.W�LQ�}5��z�lU���eqU^���B���zA�9#Y��g�����k0G�q����P!{'&�.��%����^�W�ۃ'�Q�\��y0�O���a�M�r��F�s�v��D�<�~@4d��H��ʠ���$�t&��P͠�\��<
o��̧˃[k�,�pͻ��DSO��Z3ɟBW�{�J�M����l�56o�h�:����h������0�=��\��U������"K�vpt�i���
��o7��N�Q*D����$�����U��f�G^4����#� �'��� R���Dµ��x�P q�ôL'�]':��RB��CF8He��|����@`/MS��e��[J锱	kP�)�N��2�^�ݲ��D�� %���De�ϞFn�]Ϩ|h2�ֹ�7#��O��uh����Y}��ƟZ��ğ)۝&9!�.F�v$2۷������dZaR�����he�ZD׽B��|_���U�_�$j��z앾�W��s�F���b�Mρ���.�lmXT��ޜ�9�߻�`��w��=E��ј.�8�sӫߗ��t����;@K�I�`u��W���S�����f8+��aNq���D����|��l3����%+��!�W4����a���h������l�]u�uӴ�%Ee �N�Oі$�^&?�s�JxRB���
��锤 ��q���Q녟�|]Dx�)@�GhD⛺t��mO<��
�)x�^�T5�}jd� x�\fD/?�����k�
l P��'������<u��ih*�R�ksh6%�IJ��A�8��x?�����z92�N�7�1�y2:_��RRX�ɇ+f�)��,�,��e�������O	!�XΖ�Ң��\�s��&�8�%�>Pl���:Ψ �3�N
��ӧ��]R�?tV�`�q!w�B�̿���>fcʳ�ժ1����[E\��6B6S~�=�3r�o?�����u��F��-��9{&mA؁�_�F�`��� '鞖�X�<��i�;`IH��eD�'�8 �'�r��h(N��?���~�xO�� �b�� $s������u2�S�9���!�}��ˮ{�uj��U�R0~��-�ts��&^	@$�X6�X��1�K�9�Ç�֩�wK����H�7��lS6�J�n�vV��0�\�F�H��i(�ߞ�INi�|�O�׏�_�՝tG�HD�k�U��N¨�S ���Χ!9�b�*�/�d��\Dﷶ��*��8������DB(fs���#��&s=��s�W�h�ğs��u���k��kf�ͫ ȣ6�#"
x� r�
GC2�ۋ"��g���k��h)�ZN7���'2�;=�u��M�ۖ�_aȄ�`�SIo�dD�nB�Y����4��t��Sl���ڀ.��rx�j����9Dy%�8�*�JHJ�E�[9��f�Ğ�<:�RWo͟��B�Tv��S	ts&��QA�f�$�����m�������Ky7r�?4t�bD�֕��)�6yA��n�J]���?��L��և���@]�PLY(�<�o�l7���_�c�8ג��sZ��ϋ�L5 �o%*}�H�6�o��=�p��g��(f�NH��jk��6W�A�c=la���)��q
H�dT^����r�};��V�����+M�hZ���p���ъ�͢.uzW�k��xW���uQ��u�~���`�@9KVk}-Qn�x���89A;�5��XL^�2p�3��śM��I����P�v3�l���e���1~;"zd?�Z�9�ǵ������aO��\ ;�2 �q��R���?S�� d�؍3'l�E��}���-X+�`!�AO(g���=I���@0_h��а�I�YT���6��2�So�S�ԅ�׋q[.Od�(�$`�0o
7O��f�{�d���֭H�:.Y�Q��U7MQW#0��p4G�6D�.C$����I���1�^2)�'S�����h��q�pB�˯�i׀��dfZp�}=v2���
_z������[�k�oύ%Kˣ1�TB?�C��$�ѽKm�:}à?D�'�m`�V��(�7&�'���;��I�yq�d��0-�s��Q�Λ�'��7�va�����:���2�E�L�Ǫ��K�(`�_��y���>1��8�;A�ۅ%�/p��
��n��1�&�4!�a$j)��X��q@�h�뮇�ػ�]���V�<�� �a�w4烒g�<�c��e�$)���X���$o�~�@�@��)nZ?u�|����Pʁ�ğ��	���ʤ�=�&~S[E�ۧ���x� �"���4��ӗc���XNE�)a��e%w;���Seq��{y,'��1� 3�����,���h)F.�z.�X�q�,�}k���t�m�ڂy�+�s?iZCŦ,T���o��!"I[Y�38P^�O��P)�E�QoF�G�R+��K�,���FG����c�����3�QV\�
`I���e.�}�ރٱ�JEg�mȸ�*%o�߰��l�xq��+��⁬
�Ss��'�v��Զy�჌�`��\��L�� I��@�5���}Xm^E?�H5�L�QN��4V���޹5����Ȫ{]��B��X��������ق'T��	��|3��T��n5�G��gL����i�vfG��5��xJ�GW�A��m�����-\��:�%"	YT�;��0����ܫ<�^wR�3�βW��t�C"k#�w�}�u%d!_-It�^vV���:��c����>�Uf�j�X3��Y�>u=�ZZ˼?������9��Ӓ������}��'�F4qw`�'t��P�nی�BQ�T��Ȍ�
����W��x?�U�0G�U�b�ʲ6aȐ֯��Vs�g�}r�ڝ&�W+r�P[��1�h�IK��H�9�?�rI۽�f�hJ+�	����מ����'�}/�R#�x���=�6�,�'��BZ�E�%r�h�c �6�Xs�e�����`tAZ��?S,$�Դ;��ǶV$����&8V�Qږ�E"�ͧ�]��_j ,KED.���-%L���!����3����׀�~�ۢ�ߝ5��OJ���P4w��l�'��f��o��σ��$�{N�/�ċ����)6��d�l��ª]H�90�-��pd�=]��F��Vq�g8$�$QF�M�:q�������pr�8X�:�n�n@�)g1�E��W�j.l�)��x���O�, �k�~��,Y�O� �O�q�x��o�6�RNO��g��߃�j1Tf5]����P�~�_;��}΄/�Z���-?��oV�V�4�2��8����p�4���ӛr�x�,E���Bߋ�bE!�ȸ�n_�?�O�]`憒��k��Q��I��(su]��ү��o��n��H#�!/X4�V�+��V*H��_^�:���쪠���E��ǿT��ݰ��[j7pwT�׌���t�f<����Z	M㶥��v��J���
v���<��I��t�0��ԾU�zn;|��,��@�$I�}��B�MQ)`[T21�X�����z��4ѕ��q� J���=�wf�#�{x~���N;�Ny<6'����-]�f���x2���?���Uw��A��E�3W6�kv2/R��^Є'&,#y�*�[�#�ҝ\�-�T�nl=qw��/9lj@������Ѩ����#�Z/Z7��QgںWۥ�/����Vq�Ρx L����D���Q`��J��/�V������j]3.&��Cr;�Qp��׭� h�F9�@$�̝�U�i,��Z�*��1�$H���b')�%;}o�/u5×Q� �)!�N8ڕ�Gf�ҙc0CZQ���a�0���M�U��{���1&���`-��?(\p�	z�2P?U="L�[m�ý>wsr���ܾ �����GoK�����A� B�����K�r}(�M=��>�3��?�Q˫X�~{c$%�,���L?�؃�:��h�+���e���6���.��p�����->@�iM�i1�+��o�i�� �8&¿���7�-}����eN�8�N��ї�iJ �� ������r�%b$��ۜ�Wn�B>8V��,\>9'k�(-������}��Tnލ_2��?�>�I-a��ȵ����U���(T@�%�G����q<�(B"Hg�-�g�G|�5�����V���K:#޽���2��p��J�m�$(���J�|'
B�@��uha9�"x��� ��o�2H��U�4��{����8}ȋʸ���M&㼯0X����-�w�Z,u%-�We�*�p�.N�qR4�X�k�Gs�+��}�cbyT��+7QwM�|��>��GZI9���Uؗ�-�:�����/��L��#��
�R�kl4�jK܉�áĭK�^઀`M,kz�3����d�J�+b�����/���,�������e�w�� .�����4݁�1�P��CO]�-G��� �PW�ˠϠ�d�I)@�vih0���u�15&���9�@�#QG$ji�m)�=��P͈��;l��uD��0l9j=kZ3&9�V5�r���y��	�t��*� Gct���$5�y�"��&\��Ib���Ȓ�۬D��E3F;�^��>!��.s�M�H,J�	��9^��Ƀ�4��pwJ`���A�|o3��|�c1�}rţ����������:�i:��΍��y�/Xw�1�$���̱���[F�<|�fM VQ��(���0��:p��oɓ��F�����[�%��]'��A�E���a�R7�cc����ʼ�b^�5��O�-��t�f�-�׀>L��r�\�6b�k����h:��v��)���7=�Z6\Q�,��UN3�����t�\܌ ����%��w2�@����$<'x�~e�xL��-d��eMnV�`��=ِTT������bYR����}�J G���h�WO�J1�����CZA�,G�vn=��[8��@\����QXj�9{�������Ueg��u����z
��j����ű�oRJ�����7�{�&gS�Ѐ��Β҈�a���:Ի=ֺ����
��O�=�s�o�d\R���a� 
����$pl�ݨa
|�P˖���=$8W�9/� |�2^-��N��I�߃V�v(����FW� �P6��]�cR���mʹkϣ�n���Cd�&�xn�9h.d"hv��Yk3nl�mO��yp�p����e=�P'�$:���5����T���R�\��)5���Z��`pk��HR\�@V4luͽ��mF�Mc�P,븎7���k�����=���VR���O�S��W��⯇;���6#qq�$�8��5��q;c�1��b'6r�P���js;��. �\|<�W�\j,��o��M�^�R���/ӂ�k'&��&1V�r\�3c�o��|6L1���Xٜpv �_��(�	��۬;u�d��Z�[.^	*�Ǌ��A�+<4PFlE	Y�m<���3��OL�����ￜ+��,xP�X~�8a{�ԁ���mR;o�I-x����l�ߢM�Tgў�����ss�$|-��Ȃ�ۗ��_�(����*��3�w�dB��V3�o�1K�P�U�M��U1�6�퐢�G�Z���e�K�� mqC��O�G��u�\4[p��E�~�a�)����T?܅C�r�at�ªxm����D
w-��lh�T��KYK�V��-���vd .@*s��{��:��xG��E#��^�p ��G��`)�Y0���o���r��D�%�ݏ�?�2� �eL�7��Ĕ��p6�����Z��wM��Ǝ��</��ĈN�U��y8�����ۘ�O��SF��[�8X�����?I!���8UJ��B�<�����UݸZ�]�nsm��y']3�0F)��.^N���>-�D����iU�֬5@A����06�H�
��F�0�e��	���}U�,H��!��g�C�Cb
ƙ��� -44] ;�Dŗ�ª����_�܋i�-+�S�?���ǂ������ݠ�&=."(S�|9؞�_�aΪ ��O��~�3ըJ�A2n���W
��,��/�J���:��ǰ�1����m���Dz90�P�Aƈ{��Gl4o�/ӷ�0�x6���(@?�k@Qf���N@��1ݽ�@ГJ3����e`$R���g(^��a��,+��G�{��p)�C�Mr����Z�Վ�롮 �|��fd�����$�N�AG2S�HǬ�p�����/��]������3�|2�k�O?���xl��G�Iڂ�K�-��"sZe���_�/�X)���%Qݵ�����d�`cy�زjQ(�6-2�R��G�}n{e�t�+���A�.*j��>u�R�k�#�}��%Jr��χ��PCM>�顲�g4&��ξ*��,��:kGҀo�f�0/� vLh�� �G��oh�8w`d�ypYE,�\�/ϰ�<��V���`��'�@�쓵�/���\���!��j=wMC1��M�'����0�!m��~A�����G�-�ߑ�u�/B���Y�)j�F�s�|��=�\l�{���A;w���)�����W�������ȁ�B�� s�%�Z�o��)�;P�%��R�k����V��oi%��+p�q~�Rje����j|tt�2h}l��]��2òs9�M����?xU0�ŹȂɘ=�ssQ�̮�|iu6B�붺�Uύ'�/R	�wZ>�}�x��l2�6�́WREG���N���z�x9����y���?g�$סl�j�@���-^�sF��g�x�A;��R"��? �s���δi�*����dj�rw�}+B�}���;�i=l#˶Ȼྥ-
2��
Bӛ�6#<���0���ȏ�دe��$ �_JB!fZ<��}�Z�|�^6ݯ#��\�6�R
��o~��+�O�\$�'�^����MY��� ׃cU"ZJ�l�N�[G��fo�NrD���_]Ż��	�ܲ�h��p�����×�R< ���WcFɏT���{�Q)���a;�;%+��.*��z%�x/U��v,�.Yuc�����o�}����F�\�LbΰG��
��V��Le^�dX�@|*���d:)��,y�H�!�F��Ԋ<��PQhx�I���>�r�]���@�΂�������ʛ�KL�DF���܋�����x�}��Va4��H��'��mF����V���֕�㩈��-T}���S���Q)���H�9�}��p{N��$!��X��=B����4���NM5���{�$[';!�\Q�U�_�oP�X=�LY�@�<���<@�5�:2�m�E} 	�VFR����EРh7l�CS�zm�sk(�9��W!g�%dsY��y�Y��8?0��b<cO1jJ�`$��ڢ�c���gO�CJ5�|3Zr,�����y�g���?�3j��Oj���"��t:�V�]
�)�J{��u��<��9�9���/�����w���,��)�t79��ŞՆ�<c��x]1ݍ�������Re�-�|��z�D�������l��Ō,��~7nd��\F) ����ٔM�|*��&���/���-?[�Ĳ�X�r�}3�Ȅ$ ����a
���2�_�6�W�*b���o[��-����f[��}f�������qȪlL��Z�'/�S��ӌ{=�z_!���Gݞ�3u���ĉ�4&�0ǣ{޻�՜IcmRͷ;���$8��[*��� �!C�,��!��e����`v�}�})�:�:���crBY�u��;���ȏ J�V�aLɱ�C�!Qӎ��x�*᫧6jq�8x�+�0R�ضu�1p��~i%a`�-�L?�یN��y��9W���=�\�:+$�a��/&�[<�� ��g��k.�,�� ���<���`����P��W����2ŝ�F4��~Edg���;t	�D �l�q
G{�!(���~j��oǸ��l� �
���������O�K�ʎW~ �D/8JH�q`���)��0�ñ���Jw<�4,b�F�n�9*O�"��m3�;��q�V�c�5��cx�[s�	|�I��:�7�:��[����vTU���(U�K��B)��,�������5�������ә�a�DZ��*#ٷq�+��1ܐ�:���t�X}������\�}��ct�NW]����j�4�)} y_{���3I���g�(BP����s��W�z��{gs��\.�~�L玀����[�B㩁�q,�Cҷ��w�@'w�1$Xf#U1M�͎�m5��cx|$_���l"�Z��hE��+�a��OT!QW�����v�4��A�1�j���L��2�hw/.ݍٚ&:���:FekȲg�C�����%��V������5������A�=�]A���b��l9{���+T4	�y�R?"죹ז(�o�E��XC��˯�V ��u�Z�@CȆ�ٿ3��q�q�yͤ��gh���<!������>ՙ���FX43�ٛ�N^�� �;�XJJ�>{�{7`^_#��	��W�cZ0H4� s�&	0z���c׌�Z�m��}q��]O�M��_H���q���_஺r;��5��Ԓ15�֣�͐Sl��j_M?��g�>�i�BX�����+$�Ӏ:�ߣ=a>&�,�Cw��%�7��Ӈ�.�m���^� ��qT�wa��_��{���8>�ё T��!F��B��!�GL�<��a(�:��-�f�n�"�۠�Cr�sw����_�ɽ�H�T�荵�r<��êh�5�[����I���nު��R*O��䔅�'�|�gVj�_+V���́��.���'��}�q^$�.��S0i�PyD����\��f8ꂶ�}ʺ�`<�����I�|OB��i�.Z��v��P>,���@%�|��)8��r��2I��N:�Q�s�qU�W�	���6�9e���N�z2X'�����xU�e����X���J����?�i�@��U9�4o���S{A��2���%��R1���.*/Wݸ��Z��u�\Mvm�$BIX�2��)+����H,M����+��d�W}�4�f=��w]��"��w2�߷W���6���.%qY�)H��H$EI��zZ>!	�/���8+7/�M��C8
���m�k/�E]��-�m�6Z_鋫�8a�v��^���"���un���Z����f��4jt��/$��xR��(�7MeV��R�u�$2�y˞f�7�b�83�WUA"yg��af������{�F��>򶉊W$�qGǖ��B���Rz jqH�Iy@���ʆ|HU�=�-M�Q��3�߄	�b�ig甽�ͺ�7���{��ϼK�1!��?1�E�߱P
u-�����M}B�,:�;�,��An���|�ꆣ��*%ͽ��]��1���)hA~'^lࠋ���(j"���­%��ɏ)>����<[<XG)���l��dR)�����v_K�f�Qu�9�w�2Ӵ����8/ͨ��>��68����k��zR^��V�PPu� �9�d#}��i�;S�}��}qt�*D~x�^��hd��،�����Kr+�pM���kE�C���}6���&m���>#-��A���!8�k<����7v�Mv�ϔ�-�F�ك粱$�����&����tXm�5Ņdv	�'�tmw:�<޴ڈ!��>��pp��H�x�{/-g�V3!y��3��f"�s�V�(Wq;P���ۻc43NW5^�S�#k2��o��1��������F�K�f�>���i����q��u/�ֆ�$��2zV]�@�.	��:�D	�Rh��Ǩ�S��Mڀ�웹s�N�oAۇb�j�[��������0�#�^�7D��b:"�������{��v<^�o\?_���H�~r�zI۱��.�_�7֭�k@����4���A#	x�������8�?����,���w������_�?�ݥ�GQM%)��9*9�f�P�#Q?`w�����w�O�8v��B�l�9�O(�M����Bb<aEhK�H��
ҏ�K�O�,�h���8�U��J�[J�������<l�-/��I�&ˁc��n���P2���ܒi@ԡ9b'c��G�e�9����F��͕d�|Cn'2* r�6���_��Au��EL�F���ք����e�s?�ǣ�s�����:��l��+�h���>o{�hx(Fx6�!�FQ(K�Vc�O
r��qSǶ�.3�7i�K��Y�h��'�~����]!F��\ìu��dp�r�Yt�����1WGE ��������w�Z���VCW$��i7/�N��sio��67�D�L{l�A��9$(��,��S�H��Pi��Ǭ���qӉ��Y����
(P@K?�u%�+<z�y��N��<;�.��>�av�)��L�}ߧhH�e@��|(�]�H�?�Rb�Ts��Mpd�}���+v�y�j%�u��yo�b���sg���*5!�B�	��܍��C��k�Qˀ����Rd�l���؛��B�}��-j�/�g<?*J����9$�6'#�_:�*��"r��r*�I�U�U8�CN��le}��ª�j D[~޼��%�VR�-]��rf$U^t$�6e��ă96�^�E�-��L`�7G��򑨙�1�B�ʡ�y��zSf��2��N]~"FB
tR>�[�^��(���}�D�ל�� �v���Vm e�َ����N�r���O[\Ms��Z�b��X�}�(���!DoƝ���a�˿�J:\$�ڗu����GՏ��ǰ���K�-x�X��	�ctA���L�cHG���_���{�g��K}�A}��Gv�]���s^p=$� :��S��1Z�T;b0
k���D�_��Y򋽜�^��9�^���T���=�����
C6TܩX%�שRY�Z����7�A�c@���y�,N3�ۦ2O�����������FS~M�U3%'�i=�C�%`7w��鰶���@\��ߏAf�ݍ#������و`>h�-֌Ф�¾ Y��x㰷�^�Ch�1��Z/
Duv� Rɵ�i��H-��뒹�N�uC%������\4e"G�\E���1��{��@�L�aUF�#,�Oc�_!��v����_S!6Ɗ�Ձ��S][uN����v%+
.7d��r��di�Rw=�%�e��gN���>O�X�҃.��``��n���r��9��H�(ǵi�[��u�yˡTr����)h�Ds}y�)o:g1�(g�b^#�M�ɟJ��}߇���27�#�����|/{�Z���8xܘ����˃2!�¹.'�j��L�<�RK�q��W\��3��5i@����.a�,�#�$Y7o��2'hC��o��w،�
YZ��Y ���"�!�I�P5�:
ꅊ=t��H����Dl8��1�V�\L��|�vPpv��?1�x�&mB�����@*�-Ӄ�]$�lH����Wo�� Q�� ˩��q���Ϗb�+���c�e��%�+���[��5�e�eN�R�3Y�dS�u����^,�^�VuiM�"HIZ1�	?5�PZ���Z{�>��f�p��p!J(�p�(����>WQ${���t$G��X{��M�c��t0BB�y]�UB�ζ(V�ئWS�ơȿU�΂�U��-F�"��2�{���;�`rd� ��%JwQ.��֚�$j���K�(<6�}��U(����%J�(`�|� ������dΆ����Q|Y/��=V�aFB���x]Y�'��VpqKD�Q���R��� �wj��1!8���S��||XM�`C�%�fۃO�S��p<��)�5�Lj�J�TLw�մ���VJ6A�<W�+l�{���}���׶@�K�s�WW�z�}�G��P� ?G�@�lT�k����J=O{� �%��[�(�_o#ȜIpf�Cجo���PW|ؗ����q�c4-n��ګ7f�'�Y�x�K�X�����X}��cM�U`�Ȑ\���p* ؃��ÛE��^�)�7�5{�P�������Y���{�pP�J��ܶ4a����5Uj��R������Z��S?B%���t���@�JAⓠ�e�{�Q�0�wrOt>��.����#��Rji'>^�2��8�!�*J��<��i7d��z~YP+���[~�	��H��|����g��K�@<��+HL��a�=,NM�K�G�������I�z�椵��.{ �*;���J������V_v����NQ� ���@��������dڽ2�-D^��|\��B�S��6Q��Tt �j�A6m���F`�r�^DY�r#�L��^��X�J~�WJr�p�a %��o&o�k�o�����nr����T/�A?c\4F"��fK FU�H�A<md�dG0��{��،+��
q~� ��Og.!\%p�Ɵ]��Ѐx������S	�e�/�#Ĭe��vӷ5{�C�Y��q8���i{�ܗ�QLn����z;V�2o"<����OD��-KG�8���2Q�4JU�2:a�ϏR!�����8��-�c�Y?y��t�	"����h�=����@73��H^E�� 㐁�c�����})��C{M�'�,팽��<�SES6���ZH"��������]��z�crK�%��қ�A�M����s�2��/�ax���c��Yc`�w��A��w;(�u?_8�޵���++'Ź,�t�"9�(������d�hSΰm�D�J����@���b�.A�0`���|a�xZ8!I����5�p�7X��mp���B�����chU�8S��
�e+IĀ�����r#G?�r�;�ύ��
W�C���fq:b>���ῷ��Z�7��ͅ_g	6��5x=^߿œ�,z�^�Tu��r��!�~a�9�wV���~tQ��Z	*^��]�e�j��9�s�޳0z>���C]6�+%=K�k����鍰�fB?��u�_��/�I��`�M���	�1?1?*���י���qb<}�z���b����@��&H.Ⴑ�{���> �m�p���R��xj����cY  AV!^��8��Rt�\7���(yo��I#a�P/'��Y)UuEZ�砋م?c��-�Tm�L��.�ͤP!�=�"�8�;����c�3UZ�O�����C��8)��pB��:=z��z���)�,���V!�zw��-5x���طLwux�÷謸���,�N��A���e�t(!����,�{�_�C|Pf矋F�� �d8�D�q�m�?k��[q�f��'�7���3\�;��[^�������S�3���v�4H��*�koU���A�ǋ �N|�r&�-Y(W����5�J�Ln��X0��y� EFt�45b����#^ŝ�p�t8}G���]�
y����v/Y��v�e���
�s�#e�m36#T�A���.s��}0܊"U�u&`���qn���!h;oժ�B�To�5�{pbA?�+q��N�a��-�m��,<�sT"�ġ���f~N�rO��^x�[~D>^V��?��ɴ�(;�P
n��o���,[�Jl��\�����(ZW��.�n���}�yD�`z��w:�b~)��@��y���.�|�0�eF�6d"3�8:���I�
�@Y��ZP��ȇ9J�&X^)Z)�����(������	����q�����J��~o(��̺а~P�<Ղ�P���;�M!��jY=nC�?th���B5��� 5TJl54г1��{�1)]��Rn�$�N�*.��0}G�.�s�[�`�Y�z�)��U	+��w<�'�{,+_��-�����y~�D<�����S����0�ǄAjу���O�u���
l�<�Q�{��0T	5g��o�E�0A��`���l��Wˆ�~��8&�*"��j��zUi�[Z�Z����v�Bɴ�9�-ct�'������T{��=�����0��2tϥ�#4�����ds�1�� ���fz�!S�ߖ�ɢ��>�0���at�"g|aꅂ��ސN�l�Ǘ���ҥ.���D{�0x�	5�/�H�Ǫ-�I��e�u�x�^�p�_{:C��XZ�� C�8�2#�?�ɣQ��D�V3��I���)$2�hL<-�T3	��Q�3�����JN4֨	<����N:���	.w_q"���2�),ѳ���yD�V$r���Y�R���Լ>"����&Gr]�Q:�2bR$�^+��6Ol�k���J�}ᤷ;zU�(1m�s�u�(�|,�I�����ݰ���|�G�;\dH��������W�R��3R�����u��Y9���Ɂ�Se��
�����񣦣'u�q�}_ț�w6�O�D�PWx����)�,A{C��T� D��r.棇��7��4/�FIlw�8ߝ-�����=�WYM�ς�<�A՟�����l�6�'� ��bW@�H;=o&���w�< )l�˘;5b��fDI�p��J�S~K\o����k��=�/��lL��v$l��g�W/b�JO��2�X�ML ��g6��Fkc���o4I�ʞb9嚱Ǩ^���W]���9z�NCW�{��+$����t�N��2/)zy��lv��S�g��|��V����bZm�(�5�����<����!��DX��G
�wur�@�D��
�
��[�j��My'���	��H�]w�j/�HE�a��-�墱�W��
�&�<X䧚~D��y���l�R�Ќo
�����e\WZ|�����w�l7iZ��j�\8�6�7m|��2J��J��a~�<x�l�#Հ0��$���2��p���>b՛IB�b($��/s��΁ͻ&�3��p� �y~ȺᘇO��J-�}@�bπq����&7v��{��@�ʖ��Z�$��A�aw=��qWx�[��Ɲ(�L�	A$���j<�U��y ���&q������I}��C�	��y=���b�&��j��O�&���^���K����J@�����N>��s��'�H~��˛�ꓐx��H{�:,iuμ�h��u\��K�yL��|���͒zg[���M2��屩�/����b�_\�������甸'q]5����:"f��آ�L�m��y��L��h���[}��Gj[.�,�Js8���_;FN�>��1Svu.���j��r�>�d��(�]���3N����f����8�YTC�0o���Pn�����I�*?#�q�K6\X�?�y@�����5�I�s�o�K�mǱ�3�0q�ԍ�F�l���B�M��X��V�rP�M���׷Q,5�8}�/���>y��0i��VFs�+^ZjqQpτ>�?��<�5�0��ͥ7b���~yIXד��L���%S*�����w���jn�T1|uD[�0�X8R�#�5B��V{��'蔮�u��/��6�X���WA�U��G�6}-D�2��	­��'�3��y�������^�F�m����Z��"�Zw�pq��ZT͕DO�	�`T�}H-5ĳIɹ���*�<'�VA��`*+̩?��@����3F���]id)��1��ͼ����x����Ƞ��l�5�����wN�R0uf�
1�����p��:��Q��Jʇ�����v�&�w��nJ��� � 6�u[ �I9�>w��LFN�}&-o�V�D�KݠQ8�3t(w�j��|�)B !^�D�~ .���Eڵ��L�$����0j^�)�/,2����ڏ��� ��g6?	�ɐh��x�3�t�]�F�s㎫�}Ԯ^�*9�g�䈗1f�#E�l����#��ٙ�Ǳ�A��C4���^���u5uV=��}���\j��l�]f�Ե��H�OT��x�=�������	ȸ�u�k�+������rs�ZgF��;6�^�C��n�@�e{����O)�+��_�Z�>�1Di��eU����YYS;_b��n
0�=h/�q���6̓{��#��{43��ᒧL^,�@Q�'f�D���n���x��n�&c{y6�Ѯ(�ڢ����U���d����������¶�V�԰lw��_b�M���-M���5,��S	M^�,#>똕� ��
��5u�����a�j���1�Y��5��ۚ}3A <�w�/9C6���a��ZZ�\,B@]g�b�П��[$�$޻jU3	R�;���<(���k�����Zjv�Z��"4j2�����l��Be�w��hS�P0�bB�@��}.cB�޷��r���̪V�v�ۯe��:���T/|�4a���n��nU��'�q"�s0xl�B�k)��O�X��-!�C�(Z��a�g�|XRLQ~�q0)04?�hm2l6��)��V���@i�Iw5M�#V=�M�����W�c�������Vک�A~7�z 4H�<;� ��J��	����ʷ���ɲZ4l�,��kOF���~�,m6������{��[<��XٖH���=��at�8��m�%��B��\�S~#�_>X�?����{{�x�M�'�5,��4�Q�u�����p�,3H&Q�Tp�T�O�5�N�9�/#�"&^���-�o?+�V���JP��
�F�w�w&}��Q�D�(�w������. �?�7E�/)b�ManM*���˯a�	N��#�u���Գa�s2��"���.np��(  �����
��ֱ�����5��
+8ަ�Ԝ��a�R�	�1�x�A�X�tp�,�����Z���ɡW�N��kɦ�p'�`3�����"�@������l�i�EDذ�Őh��B
���K8AQ̡�e�_]����9H��ᱷ�η�R|!V�&�5x���Ts�t_�of6!���MqO�=�P�y����J:qMT����?®?O�s?�+��7Y;Ig��O��p�*����d�|�h�A4U�[4��2���S���_1�8 �C�~r��"��,ǽ��;���=���.��t���:]_򭴘0����o�ړcL|�&���fO�ߌ-�'�(?O�;EX�o��� ���p;@둉)��"y���
{�R�'�zb��x/������t�I����dT�I���v#0I�x�z�ls�Ѡ����xC<�����_�61sAy������W�i�%tE�룻�嵣���t ,	�� 6�"� ��%�q�R���|�hu?n9��v8;��@�d��)R\�������:�O=�t؇���2������WK�5\l������<��W��"�����E/�pK��/�F�w�p�L6v�R��z�%�C�g~�}����i��̤��-/0�T�4gL�9a���y"��z���%`z�S+��{/ �]㱂5���maď��7k`��̧������B3r[�|S��g�%�(��Ց����S�#e�Rr��g�>��]'��'�{�q�|�u��̯���3�^%�Z�}q�U�Q _p+����;�c�a��6.�cL�|�*&r� ��9�����ڃřqG$L����6B�o���6�?�-�z�Z���z؂#�S{�����A�-�:��
^˼��q{��o:_�V��H�|O�۷� �ӟ�@,�B��>i%{4���;���̶�z L�T�������x� ��
�礫J�ԟM��o4����v�l~�7@C{FvE�Fk���7װ�ތ��)g+ل�3H���T@�DK������c0-�7DV�������Z��Y��ɿ�?qz�]I0��<
�j,H띸����	YnF6�xY���E�dcBcA4��,����{c���e�.�X�*�*�;r��1�q��R�G�KU������ ���8���<��K�C�0f�C`Ë 1�B�<.�k���T�fF�&��8��1��\ڕ�{)�cg�G{��cI4��&���Q"�߆s�l��|&	��5�F!9�ӌ��o�ن<lK�|�Q.�t���U�P,Rӏ����u�l.�Gb�ݕ�i��H��XI;�9�u�1j�9�~Sz�bKV�׼BTR�E	�z����<�̓创K�~%+	<�U2�3�?������s s��+C�à�ӂf=z^��B��"�#`�=BLD��<���_;B�Fг���7��$�U�8����鮜i���_�a�D�S|u��q�ѦЏ��^�:F��tFb(+�Hd�@��C�,���$?>(�.�!�5|꒟c9���j���D��|��b�o���u���.���6$1}��I�ƈ��LHA'&�xO(����y�a����#р�K�?��x�������Z��	��M�c�#|�n�*�� ��%݀]*)���p�8���������2&R�r�@hs�Q��<����q�6,��	�����bQ0!FF�l�I��O�M9
c�	�5�	f%���z��8ߊ��vy��#��T4/#�������y��|s�/�ÿkH
�G�1�Ig���RE;Ә��n�#Q4���ذ"q�?��C;d�
Ы���|����<l�R}�E.~�_[��tD@����\Ǩ���?a<J��;+~���'χDf��	ϱ�g�5e<x`�f(�K��ǋ=����CKm���;!�)�&/�V��^��*h!%�Ũmz��o�Ӵ�d��k��/����z�A<�pweZ�MvVp!6دk����6\6Z�z�$�(h�<^?]܌����.�:$��o�Е�0���ځFV:`��œ��W=�d%�7p�.���˻W�N`�3$��_	@���qa
�W3ˌx�:��-9�w���������,:ɒ��2|]-g��h�<'��d����?��kJ�e
"c�M� ��\PТr�䯠��r�k��߄K���xS���%DیN\봇�o ��-����O���66�~Xڂ���C����x��W/[�!J���"3kh�0�M�#g����G,8�x.^���:e��>3���tTll+;���[h�1u~:�fNu�by!/��u��J�YQ�\;�Ʀ���|�/?�|j�l�y�`ֽϬ=O[_��5M���E�%��h�����.w��H���PElH�
���%���z���:>?/�Ml�]LUo��I3b�`'~���?a]W��Ԉ�P�M°莽JyW!�k�\�j�)Q�cx�v��k ��=�'��$�n�n������:������D
6;zE��t����_��D���X��g�x�vFaJ
��}f��u��[�R!	�Jh�n�q�)�1�S�_fX�z�`�d&�.r�r�i�8K6����;�@������>����3����;;G�t`o�r(q����7�y|�8�vT��2������	dYEm�8msѥ���cl�p�zk1�tW֭^8	�G�$�h�Y`b�U~A���*����������m�������:H�5m�G�Debp��#�Pw3�a�i̬���2��j_���}��_�qg��?����O��(�a4�e��'T�h<Qe���S=��:�3�� i�p�M�`#0�B^ۑ�Ը��k�}/J�d0��	���[��&1\�q*Z=�#��7��C����qлu�O~|2dE��*}a��<��\�\�ٖ#~�r'��4���pjB�p~[�i��p8�y���CrB�4Q����k������k���f�����e����������A���P�c�׊\���o$IfŃZU>xpS�4D�>�oM��m.�����g���k<�Q��<=Ɵ��¬t�Z��&m0��#�`���5���ƧUUϣ�i\B^���������6�fW����E�ޱ��_g�-�7�Hf��v(�A(�U�~iߧ�F[��ɣ�:��R� � �q�p#yml�h����gvN�gZ^���'s�(L<^a��b_اd	�7v>ik�`�r
i�� IQ�V#.؆�|�6]��ǥ�bs8��+=jp6[n7C��W�6uo���d:yF���@��[12<�Z�vm�*`2��G =�� ~�H�FU7_UQ̐����e�|��B�}0�o��u2��Ć��i�p�7m���C~�~�K����{�N��)� �C694Θ��/�F��E.`�ژ��ܒW�NG=0�W�+��:#�����yb}������du�ਖ��jҭ�I9��t��8*���)ɀL�����5�5�k���궢�M�=��� �r7
���%�� �E�F���������9֠%�H�7�3���zv���A���
����#tt�^�` E`��%�k��	��R��c�O3�+^h!��������A��0^p���bB��.D�OfqOQ�""0���)�B
>D^=s�ҁˡӋ������gD��n�2���X�#A	 ��T^z�x�Yd��D��|i�u;ҙ\�KfFY��i�2aje̥������i��p��v @)�H�4 |P-~	���g�4}���L]6�.��Kl�%)�/]�8�SK:�_���Q`M�U(���j���4s�`�����Lpn���A�F��>1g�q
;)c�0okE$��r͑�4���|���M�'0_ �L�.����V�$©<�Ƀ�]?�D���e�k�|��;��_��iC��Ҿ�c�-}P��@��cy��o>��M�����~ٴ&|�C��:�w}$���Sg�d��D_���<�����?>o�� 	�`e��~�nN���vA�4<o�hq@ં ��CE9�m9WkM먳a(0���gg�"썛T���8FGqh�jk�Q�F�|���Vʘ�}'�0.�S塊5+�`����J���ә�cI������-yh�7MIҚ� 3�8��<���zdr���.�PqL��J/��T?*�`?&u���V�r��	XDCZ����cf{ݵ�>k�|��g"�\X�7�����B�}��{͂"=g��i���މU�0_oNcBň"s��Z�r;���QN������A9<�:|@�ge��z4��:���M�ߣX��"�o�˵/�I�
i"����������p4�J�xsf�)�������K{f�.(�D��PYW�Ҥj��~�A���Q\Z��>դ�V�ߨŐ��& ���!����M�=�W��upC��1o3䛹�O�7h`�$��L(��l�K}"���:�D,H�,N�D��v-���]����h����!޸~�vv����.�h�K9�iEp �]�9�S:9?A��O�W+��yR�lN&�U�g�� ��xO-�wB�ݴ���Pİ�����D��A��Iّ���0
�F"K��\4��Nq�����2&7*���
��"H_�R���h�t�t]6�G���n��I�(�6 Pap��A��#� ���� �YZ���@0�Ud��w�cb�p�-���<��jr�&��o�V��֢D�i��I�<d��,����#�S�G���<_\�a9��j����ٺ�>���-2p�JSmWYs�_�cW�p���XCy4C$��۱��ZVPzջ~cw豻 j����-x� >�teS��Gb����҇B�li1C;�.hne�n��s$���;]
�e`����6�l�q\�6�i�j�JS�9LU7~E��w��K8N� ��#�����b�S�����`�'�$:Ijƨ5�s66Z��g�7�n1�z�Oh���O�T�K5�P�MmS�E�u773�A���	��uR�<��=s���)K�2j��>Q����XK��Ô�"r~�3��O4R��r����q�O�Wy��2 �cE �G���?x��F(l�%X�ek��?
��ܫ/��vL���~$T�l��n��W�|~����#xy��E���'�4L/�+ղ����'xlU| XC�pX���p
7d���?�'��Џ��"��"_�Vo�k�eHjh �C�Oeoo� �H\��U�h9�[�Y�����eR1 ��z�qa�AF�����8{�Tuky�q�Gq�+��n?�o6� �ٚ���>9+;=XY�>��cI�n�1<B�'���_i"��&��Q�A����t[�i�.u���W�k��GǓ�N,�~������PͰ�AzBi���!B�}�?b�6dy'w�lP�\�`}�LE!�� ���0�^�����i�����v�)H��IFO�%��q��mD�ߔ��8��5n2n�7�`
\�}̋�MkCcD��7�j�b�k���΂S��f?l,�fU��2��KVwq�u�p��u)�Y8!����Է�I�@�!�3܊j:m�;��i� �*˔ߋ�T��E�J=�k�f��&�꿛��o��J��A2s�����.cJń���q6|�����������\Y_s���A=���X��//#�'�&�����z醒;r�t�,�ẛ_g�K2�T��D�A��!$�:����R��4���!��_羪��I�v(����d���~|���}�^JO2A[���i9��U���������3��^�o�q>imz��E���|z��uv����C9���)T_�Ax����"ϡ%nZu�]�F�������c[�R���dW��?���ZV�X�l#�(���߱۽��"�H�уC�=Yb`�D��]>FI���6�]1�߿��t繢wݿھ���zʿp�)��͛U�L����$o�_�έ2-�.H3"���zf4!����+�	K3�K��q9��e̵�6;������[M�\��"���T��'Q��X�q'�"j��6SS};C}�|��J�K�~1y^Dʊ��/�����;o3�v��O/VY���t.�8�]�S��~�����ʭ�ET ���=�kr�ˁ}`�p�U�^Bu��poF|*���K-n<@/O�����٬��9}[���`�B<���i�I���ș%�DZ$���ɡu�kẇ%��ϴ�-�
���t���?)7�e.��/%��	�P�R�iC�ľ��WVUE�6iF!���Zy?s�2�4|<�����p�
�jD��1X�SU��EO8S��D���b'5���̘�T�8Z��������7�%�r��k����c=�2hS3�>�'.����,�!2��޿��ς�A��׿{�E_+�֭��<x[��u��k�����;'��%��iYSS�bꈅ&L�*Ky|�fyRګ�D��$��R��#�������%�ڻP)�#�֞L�XǑ�V��Y>�ӂ_Ũ���(���%�EKJ��T�h�l����R)�bK4�G����S�*Q@C��_GY��^+��R1��:��)h��w�oDX��!R?Q�5�wX)a_3�Zz�Ɠ(EHa�V!�=΃�S�C��70[�� 8QC���+�tF[+iN�+���/QI�\���Z��k�%a��>���,��yp�:>hK��wzq�n�Q�Rya��bb,�0R���A^l@�2Nl���#��N�nA�Ѭ��Do/ނ��?𝸔O3"O2���ŷ��i�i/�c�5��/G\�1�U(�5�r7&��\�^�T��;D;h�r�]RX�w�\k�G.KT�+��/�.�ɥ��(����E�5>d�)�S"�$ބ6�C@���qȫ�8 ��1��:���"/pu�'n�k�ͯ�N��y�}q]��k�{���-��mve/+�E	7�#[��vi���r磫 �m��o)@+�O��ϔ����Lbju�J�֌e@��:�9�;<26�,(r����cGf��(����8�C��r�B���V�I���ʕ�X��ڎ��pT�ɍ0�����,�s�K넉��1z��u��o��5q�� q���b��N����|0��ɝ���;�9T%Rg�C������������
�WC�겝��H�p�YC=� �g]=gN��3���]�L<�<�T>ׄ�}J�!g3���p��qL�QC��� ��^�+�K��\����g���)���a6�В4>����9�_M����>O�7����2���*�İU AO}�=�qs���+����<�r�r��� �9�%�[���8�5~&J#�N5$�4��Q���&ER�����>��6H�H�g��$JCn��Е@� �Q�^��%��"�kqيw���|�v�|�2H#	_�����2WD�{���qJ�\Zz�O���E)?S&����R���|�������#BKYpԻnO�	�E���TVZ�I;_� �Պ����2r��BH�	δ�d> ��ȭ�1{�����'²jK���UN5��s���T%����WˌE�t�e�.C�#O)�#D�T'�UQn�/�7���F���R51�+��NaCӬ��
����&�'���:$��C^�(9��)6�Y�d�'Z.�e�z2�V��]�\��L$<-�V���NhAr �4l��"�q{Ҟy�Fu�~����^���W*��~$vڕ�pC��i6�%�s�j'Q7��S-s���8����lz�����WOAQ�^IA�<��uʸA�B�ڇ�d���A���Dbx3�i-R���XM�&)4���'׋S�W�N�}w6�)�q�F�U'h܍����J���vM^߰�[]����źחi��*z�F�[3*+z�/���{��E�
؋��'���1(3�����O��  EX��}��6��d�ޱ~�hcIg�*Dы�q��X|�A����ǡ(
�xqJNA�a��j>��cnnǉ~x=�v�٥S%a������L��ͪ������$�V(��L�L<bWh�W�Z� �u�4��T��S�L�,� ,����f�6݁D�]�_s������r(ZN��9��G��|L���<�&���7$M���q;����K�Q�H�rڛ� �M����N��,P�kӡZ�ƻ���u`n�̯:8��p�ܛ�[mc��"����M%�/Ԋc���l�)\�V���eF T������|�B��B��
�X*`XΓ�I���b��������%x�	Z`~l�"U���U�d�6��-�Y��w���G���Z��6�j�6c��ɖ���M�b��Lj4��%��w
���Y?��K@��2gX��]\���a{��}xv�f���C#G�<��Y�5v꧃t��kt�E��ӿ��F��L&n�i��
7ȕ��i��5u<��/�y�H5I�G��'G2B�5�ɱ�ы�i[��@��WK��zg��@�����v����DbR)}��jC��j�����M�ݦX�,����L�ı��dq���[�ЧZ��Fv�2�_7ط�i��B]D�?篘"�<���[j�}���,�~*� �O7��nQDX�2:@��H
��㎲�h�N��s���r��;�H�}���)�Kr�*�и�3
�-v<���Tr������ї=7{�=��3�x)2]�'H�6����8�N %_��Adp!�o�;��j���:x��Q �8g���hDR�׶]D�ҩq�[v\
���#��w4�`�wy���{�K�q�Y���x[�}��b�Wޭ�[]�����~F�t�t�u^Q֧Y@��xj�[�u�5nROe�a�T-���&/�ے>��ֈ����y���<�w�[��/�tȽñ�=���9���>+
ؓg��z�@����Y�_XX��'V�0ܓ�wa[vB��w���wz+�PXRF,�����["WF��\<4JG�vR+%;�(d,\\��l�z�@J�ƌ�%)w9�`
Ӕē��0e�}(�Q� A���%��D�0�BG��+���t�+eR���2�R�QC�̕K���s��u#�2 ��D�Y�n�������E͊�I�O�h����h<8�_��qD7����A'Ƙ5f��s��F�Y�%�7�8�&�����@Vj�3l�,�����Rf���U�?��N�}�r&A=�������.Ñ#ji��],�mw�I�Uu����6a��d�X�l�a�t0����^�bkw�܅��(��#���|�4�	t` ���A�)�FΌ��#��ϟ)�z�?ᛥ
d;�1E�I gt��ݫC��`$���!����n�3z΂��E'��) ��-#��X���jBq6jE�Bk1�o�8]�6Z����O���0�6��7u3�Up������r��(�������o$<�%�`~��&4h�K�0:�N �`*����D��Vn���Sz�n����>[��P+1��osp���^62c�K���*���o��; X��֖�p��"8L�f"�6�# ��h�Ҩ6��L��y����B���F�YQk�=���ϖ���3���X���crw���T��ˌ&�$�
V�Y��J��%��>X&���/$�d��������*�Z�%ؤ<���Y(����A���<��|VL���T�����!�e���S��$���1XBs�{Q{�	�	`]b��]��N
�c�U �������G�SP4�󺔬�myy������7)�����R�	ξ�V2OW���OV�d�H�=<��f�,T�W8�4/�%��&CJ'ySc�֢ .��);Q�K����c�� ��gC%ny�/�yڨڍ�:��jx�%�e���T�M����*S����WJֽ!��~I�V\�b�*���[ݒ)��	9Z+3b��O�ii����r���W���>��ݩ�Eua�dL����èrg�����]3��2���0:P��RS��/؊w�&�\/�c���~�&a4h,�	&����ѿӼ�ޭ&�Cfpj��Y�$�[|�x �7�/ZV���G�A��&�&��LǇȭ�O����ȨB:n�= �	@=�U�)�֓�lDTZY���U��y��da��N�al�N�"���? �s.t���<��N���>���^� /�v���Ԧ�֦�=�B+ ~����Nr) �hE�9�����f��mbZI�[!nj��n&��wy��v*���94�^ R�V�IC*���Q�1�&P�ӟ����������s^��	o
��3�kF
������ʐ���v)��"���[5(�A�흦:&�����C2��O�3z`b��O�Z#�i����<iʏ���'�Q��cС�l�F��$w���v�%>�����Re�����*�F�&�ؙ2U`�� [��b/rξ,9h[�f��}� ��%�ĥŤ	���_M^��i	^�L�UĖ�O��X���f�<9Q��Q.[�d~k�ƽ����jsz�y��։̿�V-�Z?���f���Er:�O��Ϣ��K3�%��gk;0R����,p=q�&'��/��w�O���r
�e �b�/��w���⍮o�s�D�k�V���cz����]�`��KN����ifR��_Q������Uc�2w�E��Թz�3�j+Ne��k����|�����[�R���ð\B�?�0�z9W�|��� �enhq�P�^��=�{�o�$?h��K���)��7S���N|:����@���	����OB;:<�r y����J�-�\�^z����'D����l���]u&���s;1��*���&�mM�z�7#E^2��4Onv9��(���A��}A�
/O�k�4]��]h�5�����%�P�pU%Q8%j�￐�5\#����l z.�Mħ�K뭓�g���9VY���3�"��$����E���;�Nf���Ϻ���;�4eF�i3RL(�Z�Pu�9�as��Ιy� i�A��<�_�,�/'�+-Ör[�����1NҚ�D�r	��0�������\���v72e�8*�#P�σߡ���m��YB�a�ͤ֔��M�4V��dϗ%�ńY��byG	 ��J�T��kq*={��	X-�A����o��0��U�L��҉��@`0�:���_D��e���A�� ph���{�4��(!c���&��EWcI%����_��wr�������gg��I������kהz5h�q�SUw����pԉ����z:��t�Yy� &w��u4 Ѽau���Ͳpn5Br�x���S��$����;�Y����6�t��")S�%)ě�|�+k�	B�� 8rYA$G�'5� �L���� Ψ�p�
a�����̣���/0ؼ��R�������0+�Ȥ���};�%�mЁ�d8�'W�7�T`F���/�#w�n���~�W����C��-M=�J�`�Y�
RC����p�k�Fy�!����d�?��8���u�*��$�Q��:���/����cv�.t?W�1��`���DK�X;���Y�T�q�����}�K��O�eL�D��յ.L�j� 9wr����	օse��X� ))\U�V�{/��^ĸ��M?Ѧ=B�-\f���:Ψ��vԪ�x}�&i����f��Q���+�Ƅ�=w�pT+1�j�/mU��r���d端��c
�ޥ�vXޑ�)���ÎM��V2����~�jĪܜu�� �c�3h��Dbռ]��E
I���g��Kr�QK��,��oӍG[(�G.��swhZ�t�<Ky�mJ�b��"baV˝����`{�qs}�V��R?,��ob�+����W#���x	p�1�w[~e�W53	�|�Bİ�{Ic���%@��5�.:�ާ�?z�&�AK��4��hAv��"��Bb��CP���>�����sP��Q4�A�ƊG���il-���F����8Qa�اm}���>4�B�o/ş�pݚ�݈��/y^�";7���-@��%5�nQ��fW�̸~G�hO;��>�=��+��q�t�;)�/e����?���d��2�Uz�I>׷�(Z�ᾖ)��]6���eH��i�{F,]�/�Yb7X���@H!'�����<��;��`ڊ���HC�kg�%����H�7P���s�����D�[����0�M���ْ���ń0H+`@ s��=���I�M��2l{�ރ�D���|1\5���
DlK���V�0~���+4rR�{�D�	`Ê���HH�.�"��L���`��\M$}�k϶u�7����F@cSJ+���ډ���5��a��>���E��w�.�lYз���z<��6��@� �Ix�	�4����	|*�+ClVx8�E����_{5�O�$J`ʢkW�����U*�>v;tq�+;��&DHg���SW�亃�N�%�\�uL�,6���c��Β��~7��x���қ�^�-k�w�a}��í��V�>nP]g.��^����l�(ð�~�0 x��W�ڕ~����cS�(�H������[�'�suV)D�D���[�������W\S�}�"Y��X�Zvg�a���~����U�~S8�4~o�Eڞg����p��q�ҩ^.��LD�����h�����Eʛ�Q���A��sꠎ�S�B���KČ�Q1o��6|�:�~Nw�H���k����e%h�rE����?�Un�(��[@_?\��+�w�ָVb�I���eݖJf_bU�ԑ���@��&Bֹu_�c�ћ0�-��(��~���(ł�U��/ۿ�!#H���d�����S���0��y �0������}�t�j�ʃ�{VX�l����N3!��}&��n�3=��Nk���ըS7Iv�\z��B�ӈ��?�[������Y���;*�,�yo�3S���t4�����{)�Ɩ%�/�N��b�v���s��eۮ�;�V�K�so7�&n��`�WL���
k D�~�M~h�h!ٍ���g�i_ܟ9�?f��u�?w�p�Y��7�l~א�OhF!b}��a�	�w7K�ct ߎKuQ$&G����%1�i{8��T�,��P�a�a�����B+��P�����;,�dZ��g�{;�Y��s�l���>W��^[��bT��C�0��\PКǝ_��S���:Y�S���~���<�Kr�3�}7�c�{��6�[�%�0�ae�0��r�~�f���^�n�~�9]�������n��l��=���~#~;g}���ެ7���xo8!c�h���F6����3	94,�4����FA8�{�&���=�r�i��D9+�\V�]�>�o�z���A/ 2i�r��!P��M���ذ���c��D�\��:���5ψDo���J�r��h�� ̜���u�$��S� 7qPу���#�l 	���?���hǠ,��#+b<��W����]c��*�Qn�܈m� D�虩��Q��J�YD�N���60
���'�o.�NgI�Ľ�ܨ����4��f?#�O�I.T'���=�����m��?�^�%U;���|q˲�.��dĵ�٤Y��$p�������ˇ��,�{!���>���CN�?��P�hy�y���^n��0�^���D�%?BVB)�B��m���w�:�`���G�����oL��@.�r6������:^��jQ��$�\� �_��X˺{j(��z14��#���[W�E�!4���U��c��側�k�~�G=��z^6A�u\���Pim���Է�W����i���j��@"4]�����ER%j�f�A�%��d�LV �%2�]!�vWv��� �l�z�h
���k7�j�}ٍ���ҋ�i,���L�b,#����F���6a>R/R��:a�s{Ȧ}���˩`r{������\Ď��#
n�N�Nl��7N�?��7�sg����=)����	�N}�tOHج�Q����Ҭ����Z��#Y��/*$�-�]��YI�	���E$����Ln�̝΍�퉜�1ga�kTJ�b��5�J��'\� �+��Nݥ���c��A���g�@2)��]��ҭ߶�&_PV��ˎv����wk���V� �j��Bн=�K	t��Ay��D�`p�"@���զ�QO��ٽ�I�FQt{�̋L�$�V��r>�%q���"Q�}+���!��Y6p����T� �L���NSyr���s'L��ܶ�'h�C�rj���-�,\d���2������# �5���.j��"��C�|�I�'�2$_��6���K�%<<�[�)Jd]@}�e��g_�y�+��畿=���kQV���ؙ�K.�f᎚`"���5{{A�M
�^�ѽ�D��0ґ�?����w��aܼ�p�*�`?r�4(?��]�:�`�f;d1����g����3"�V�_\��Ruxd{��|q��2f#���;�^���b�rĦ���7ڧ�?�/�`tB�k��e=�z�U,�T�k��`>Ũ�o����m�<���m+0P�W��Qʺ��|�O�Y�3�`o]���׻[�{�}+j.�)�|��#�q7�R�V��Mؔqt譧E��DL��\�	�s���7�ιm;<���1��%�}���D������<يG�~!I��S�O���� ]
����K@���E�"j��K�W�|�B
em+��@ޕI�J��{%�L ���+�02��Ð��h|
�WB����!��,��N��V���3�5)�ӑ`u?h]�
�B��E��wMZA�N|�Fp��&9��,+y��޴D�q�.vH�*3�Tl ���"f���mX���W�} m���z��J4_;�6�x%ԝ�Iډ���;��E¶���=�i�#��t$us�b�v}P�[w�^QŢ(�O�2�I������Wb���߫G�Py:��	g\'r4|�],�Ƙc*�0o)Bꥬ�)!����y��O�Ñx�X�DR$`�Ԋ��'��ੈ��A��J�x�2�7�)�;�_艫/9L;P����b�]�i���Pq/Z!���$JI�f�9c
u��e�3=t�İx!�X��/wp��S6�}��2�T�d��E�
u.��	���bh� Dحf�����Eo������X!��p������\<Q�N�2��#ȏ��ѠƕZ���iz�3�3)c�� �]���&X�n�|���M �a-��U���u&�����2�`56ZU�����W�\*��k�����2D�\K	-�3>p,��͑�t�Իʟ����P�Մ�d!T>`h,�j��u�Ϛ���PQ�5�64��wb�9(��ߌO�@�&۝F�nNF�a��G�?�}+�ߘ�.V!.Z>$́gyD��A֎�0��5�m���$��PIڸ������(vRl���IJ�����K'ui���grZ�RY>CTs�RԐA.Ve �V�e
�}�*�L
`��o;��'9��34��h�=�s�i\�R����5k���7v��`�:��'��w�l���6˓v�)a���Zߝ��͵�E���^��sB�:U�,'5�3,���V=����3�B"k;�k.zz~��=��
0��T�+0�?�p,��N �u�&��1W�6�=H��;�)_p����X�*;F�������R��7��.&Vַ�c�L5�b���h��,�1�Q����f�.�xyHO�F�t(��I
���X���z���F��.�����T�`�qH>iL/����S������Յ@ե
�/>_W�t"g�5d k��]��4{2wm�S6�*�\Pa"��糶O;<��3�.�I�v&n�J����n��P�g�J�T�2���r���I4�a���Kfٽ
�_�(��l��	����NT/���m�_Ϡ)�5��2T��:6���V��Z\.�2�f��8����n(���_b0΢@6�2vn�������	�I��k�Lݵ�z��L���/��yC?�Z���k��94&Ev�|+��[J*����	b:�ϼ�q:���3fh@�����g�D�vb�T�;F,�%�E±���"Q�D�o��.6�
ڣ+�gs��2/����].��P��޸H�'t`�O���YūP�f~�G�ht���^N?��6GU��&�wޡf���<M�;V�'քfل�ǩ��Ėg�(�������8�=t���"�@*��-�b5��E Y�&����cp����>q��,U�������Z����/�>���m�Y)��#U)�g� ��� �^�H�(^+�NK�fqd������S�/�3�ET�HӎE�ѧ{�/�;ne�׿�&(���G�T� )��x.МnK+�V������'�4rx��&�1@(�i+}O�)-E
��F�A���q�Qo�*�3<}h	�a[�2^j�l5}w�I��4�i&��]����W�xG�>��,��M���$Z���<���Dv�>�Ӏ�g�.,�X�����C{�/�#PK:�/ޫ��4?�^*�' 4����,���%��%{�zu�;��g8� f�]�Y��4����L�p"�b��Ђ�eM���
��臹u�L Q�Y!?�����{VZun��Ou*��M�M���F��ͧ�f��.C.�6��6���qA���yX\�-��wN�	�뚒m,(3�<Zp�85~�)�3�U�<��IӶ��#$���)��o2�ے���Wƾ�%c�l��B@��U���j���=�(�\�"��wxD��
8},=��U�&ҹ���=)�ߺ���l;�X�N�k2w39�/��CVA7͸/3'������#%�x�6#9���~���b�=ʒ���f���l�>"�Tz5����f��K%"�:�P�7� �l���^a຀ͦÌ�UuAT���Wx�49ni]�>x!�|�P�v����Mf�*���:�Ȝ+�E� Z��W�ou@�kq���.{)����Gn���)ư�Yg׭$>%�Y���[(��x��Q��HSwŸ�>=^/���֫}�<s�;`��G��`�X�!4����E_�O�:.��ĕ���Q&�Q)���Z~�	YՕ�>���ك����]�~̘yH�./ѰN`I9���C���_�i(�����B㮅2/g��^�C#<-����6'�C懼FS]�P!��FJ�?9i%Aٟ/����>ސ��J[G����ψ?N�g��I>�d���Wn~��6y��ΐЙAm ��d�)��'��r/���M�L�x����5.�E�y6�]�Z�Zt�Ę�ط�B#�S�E�����wY/v��g���dw�7���"YcBV|��5=(swA÷n���)�ׅ���3|���ֺP�%.��S�t>^<�EĞ���Uء[�7 BW�Et��.@�h�SCT:���|�uQ�m`��DK,2���W��W��'D�;����y�%�Q��S�Mq"f�s@y'���Mjc)�@y�bv�XR=��]�N��vP`_1��[2[�5<���wJ>�A�{��owW��<��&�f�7�2�������hx��C�H�Q+���\6���G�տ����6�l�b|����DR9����b`Ϳ�ez�����V�94�b+�����즰���=���o�&��[�g�7��]�
	Z}����߳�K�\vR���y���dUD�/��z���y�dZ�*��	礣�8���O��RK�,��>{�$lAk~ܔn����8�謁��W��
։�KM���E��!.�C�BN��n#����(I��{̗(܁ ���!�I�4�2HƑ5��k�Pfzo��T�����v��v�t�&ZX�F0�VwZ;��z��ބ�5�N�-'�nKa��+���!����s�7I�n��X���-�M��-�1�35յ�Ҍ����䉨��1��3�e�g^��Y����Nd��cU)�^V�{h�4�d�!0������c�Uf��ς�M� X�-Ṃg?���f��X��bx�݌AT�u�s�����J���$��ޔ�oW����
�7{����"��O�36"�ZW^|,�-.��.BE�:YDL�2� e���2�j8�:O��0/���G��<ܺ�wBW�k�i��Qf���&��X�l��lXF �H��!,��m�)���~�az᱌*dOį���ߖ���v����˽��ե��L׿����Z�Ndrhة��;��ݫ��e����T
�50r!5�3�6T��j�4ޔ�H?��~a�&X�*ض���ߵH{���}��^��!y����H�%]�PZ�Z.��[�R�ǧ�7�����\�rb�n�6b�y���^���������-�O~����i��w�U
�HI��|9���WH��)-��å���tsӖ0d����wv�?.3R��>j:�iMw M�?��%����'gX��,������(��-�r���^Ç���~c�����*#:�,�T� �_'���o�n�_�h�*��R��^���oQ�$��o�������&#�?�'��=��߶_lh��!;�s[��˖R�ɸ1�A����Vq��O����!49�Lt�?����"�U%"����¦o��Ёu�}�5Iݔ=a9�cy���+B.��ހ/�uTR�Ha��z ��J���Ӏn1^C|sZ.�����H�DR�cPd��o;`^�uC�%�e-d��Y��
͹*v�Z�K2���w���==�ܯ��zIHd���nHш�����7�ͱ��ҷ�0~��uU��<�OՊ�(Ղ�1�zs㮹}F��u�V�`�fb��$�ǂ��csaӡ�bV��I$�9W�;�������S����4���?g3l�4"0��{ܼz3�K���X/C�;������O ���'��U�`�!28nM� �ǈ݊nw:�捴����x2ȼ�W>���3�"&P��NG��O�o�))��~����vՀ���L���E;��~�bwx�o ���b �.�ƙ�����HYP��-S���w>�$�� ��'��j.za-�rC):�i�T�uo�҄~�	�F3I1�W�T���Ag�mH6T��n���k�����$�~��f�P���5kFwW���3o�6���lbcT��x(����%��7ϐ���lܔ�dB���Hσ��s���0LgCA�~N����Q�4�.Cg������"V�����f����̱̐��������������@넎^J�B�oJ
?㻉��&Hī���R�J�v�2ڎo����<�j������F)=a�[$߄�V'����O�g��:Y�����ܬ� �e-�7�t�nVٞ�.�AB���=w$�(W�`8/���J�� �^���5r�e>(�Op��z�Wx�#g����P��LS�+�bY��A�`e�>>%�L঺��D^�a��8�mr�q��Qg�8VҬ��5��?��Q�M��tC^��ʓx8a�EKZ6q�!u�Jsۛn����~����\4�  �������OO��m�qe��N������g�3l��v�q�Q��qi��l*�U �iS���1?ٮH���gC�.�k�|{Y�[7��]�
|����C�����Y�6 ��h�dB�1�^�e�t�]1#�	Mq�V��y��/��ԃnY�2���j�7����Vv�N�O�0��S3xY����@�A0�P�F�`��O�]�@b>!Ecg<p�3�~u����e}���x��O����~��|�F�|�M��vלrl-]��Ge��tW�k��O/z�E	���ۤa
�a���x�)\L4"�r�����j���X���!�!C����YD�|�%y���k��C�����p�\�}`���R�N ��7� Vʰ��X��A�xފCǚ��n�u]�N}{���=g��o!}�����|�U����=`1�>DbY�T��YaaޯDI���1�-	�.����%Rc�]�����@^W���v���F^H@X��\�����e,��svc�}$Dc�Y����%V\"ѻ���1�w�[c�"�I>b1s�2����q���q׾�Z�Ԫo�ӌ'���-y��F��w�"����ȽL�AT�O,����O-g���f7+�ΰ.s7�"�GA�:��ϧ��v��RP�M���czul���:�\������3Z��X�����KX/�����c���D�����X*�EgN�B1��6ǲ�͈������n�E`v:tnѫ���r��%q�ͩ�_����#��hQaU&5�������Ip���϶O?^mn�)�)��'���^��SGje��sZ���H��-�n�W�XV�*���;�]���c��{+U5T_gSɦ�$�p����V�ø�&6�?�Τ��?���M"��Y�����u@�������뛌�.����	Ŝ�]��[��G����\����6T�z ���1�h)��dB&�W����a\�B�'�4`���m���f����؞L2-�>�DV�Qs�ה@�;�	hisD������#t�%���^D^f+�b��σ���hƠv���G�'�g���@_���e5�(�V!���B/���R�o��"u���{�>jL�F#&���{���(��yy�U [s�s���O��G/��4z@L{������������}��c��*��Q��A�U_Y�ً�����TdhÉP�ц�g6�Ę��Y~��K� �$ �=7�ĻT��7�.����@�@��$_Kڸh? ~D��wg���R٭�:�T����__,���AHP��]5u!�����=�c��RUfg�ɒ�� ��y4q����|�<�,�Q��3�2���.v$���6|��ë|�
Ľ��u����>�V��=�R�sA�vQȝ�Q�VbA�U�������6�K/�N�k�Op�z\��K�B��!���%b>����˔��:��(���s�%�´������VM4:���m�s3IǕDG��������<t+���K�E!�9��5�|����o\$�J6���������W��f�asdhX���]�31-�ǀSK�
�TCRM�M	=�	+L�:�؋���6�����C�h�z$�}�E�l�J�<g���^g�R]�Oւ��)�|�#Ũ�|��J�BR�:�V�=/�J����on2th�!M\��n�OV�����Z\�(����v�(C��EY���p	C@�d=u4lZ�Zg��M>��=��'�/�|�����)�TW��O�5��͵hG�X��{����O�c�����Q�>h�n��X8U�u�Y��y�,
9�ѧ���~e:��n{!D�=�����a�!I�[��}(E�(F(}b�z�.'�yxb�	=�.rU�J���k^�M�GI����m�:Ӎ?�����'*	��;�{&��*�\
�>����(�i=�V�v
�y�$����|m �٬�����w�bw�`Oowkq�v�#��iuݻ����~M�A��?%�P����W�4߿�n�����,�{�1��g�k����s����"�J
p�]7��Bn����9�Q���'��^�%�f1so�HUB(�&�lT6��$8i��Z_eI�l�
�݆r<�?GDR _��b�r=��L���\F�u�Ǵ?x�E3��
�#��s�cH�b,��h�Y?q�e��E$\j\�p�s[�h����|�:�>� �C�P�:�]y*�3ҚU�l�u����1uT'�P0̹7{6�ā�Hb_�<y8*JL����(�
�g6�b��kY�Ą�C�p��m�,��^!�W��8O���nyφVG��Ԉ �"
S���m�q�(��-�|�ޥ{�:�#��0^Rz(�x�΂�Vb��o������$�dU<фZ����
���Q̺����`F�M�A�MLR5��m���)�"6�Ai�9��:/������|�sM����"�IL���3�[��ӹ8`�J�.��t~�\�5b�W_�ĥQ�cH�讍[�Ŧ�^�m?�vɎmG������m��j{��ݣ�͆j԰�.���ޝ��ԍ4��¿��ޥ�~@�b��n\Xl�i��:�O5^� m�&B��v���<"� ̵>ۀ lu��9�6󢑿�^�"7�a۶F�m������7�/U�YA�O�x燄��/�l���ȹ�VY�dH�$�q	�O=���&��.��E%����][һ�s�jw���?#�w����V��D�ķ,Sc9�2	�׆�F�Q���ڏ��*[u���'^I){�\j"�ⶬ��"�]�����@�s�9�A>І��tm����yn�o�V�����hI/+��P�����ǭ����Uf2Kj���*�
,![��	���K,�:qz�e�0����WL�7A<�s-]�</,GFz(${-��T|���Ŝ�'u���ä��!H_>���ń,P��XR������z�����k�,�2z�*��Ƹ7{73@�"49��,H��3�v7�g�N��W\��w3NnXi �N'R�3M�<�Ri &�1��,��\�$����?�<�4�C5y���e�ĩ��2,����F�0�Vv5�p��^�!M��p?�Ɣ��N�V��3���b��8\%c���R�Z%�)�_��~-x��F���u��[=�3�(��_@gh���z�+�d1�dE��o�q��`�1��&�!Rv��G1̱.���I�9�B�(��tΌ�F��"��_�$�Tr�O��>Z)ϟB=D�6*�6��*�����HU�q����:b)kc.ay����C'E�d.7�C�־2W��!ڈ����\��?4������lk4@�c��������� 镻��~�2��=��T �������A�T�9H��6��xV#�(����s��m1;fJ�����L坍��Rƃ��@�%	����I =�5b.C!{�)v�>j�	���I�yZ1��ᣒ�
�	�6���3 � ��
��$�?0J���I���ް��P�9��^0q����7u�oMP��h�_�����kc��T[�O���%_�oRD�N��4M����t�:a�uE/�yͪKo�YkoT��.~ȶ�(w���������g�Ϊఖ����3��e�9���JԉW*[�%(�M4�}��;K�a���Y���jO�,��dETÙ⩦*�;0+�WIPT!|8Q�=�.�YX%�ah�DR8ץ�w[������.��=R��Of��z#>,�[q�,Ujz&?U�\v"T'2H'�~�f�x�]��!M,��h3\	mG@���t���YX�s�<!h�A��عm%��D˜��_��#����.L����'z��J��O3�(ְe��S$dP~��j���������U�A���>�ޝ�Y��e�tD �c�]��Е���6<��U�}���23�􇠹��n�?�[�/�R�Za7�o�|������(��E�x����j��I��z{(��G#	�Da]���Zʑ����c��4T�u�0���M�)�(��[8o�$\�.�ssݢ��X�0�$k�?���GR�&�6Q0���h��=�jO���Q�L�f�S�rK���=�X����*�:��+��yK߲�h��O�
st"�A�4��F��%:�W��-��YN��`��GD�,�i�D&k*�
���M �S b4�*�ŌVf�Ey�?��^:�0wd�*m(ܳ�d��;�'\�Ҩ�ed=<3���L([�	��ú-��$z|�ȹ���N�~�d<��|�ml	|��U#���
Xi����0Fp�����k-�7���:v��,7���MK9�ę�U���R��ܲ�� H�Diϫ�T6iR�L�H��CfE)�1���<��wFP�L�js���A!a|
tRZ�5�)� i�z���i����	��ݻ���!y�^���L��۟�����fk��Ȯ)� ��H�T�����n�A��(���k=(LdE!o2�*O��x�zs��>3�7�A�Pg�X&f ���蔪i�<u
q�m�fx)�&1�}�D�p�����V�P:E&2.J��'=�b(�����{�(�Q�μ}9q淃}�~�.e6K%z4f��<aa; �X�g�J�<��t��A���(Ře5�`S���X�w(C]��JT6�sG��M���5Ϝz����#��U)6!$&Ѿk~���^��'fO@���890�G�_/�~}(��K���<����е�kw!`��O�M�m���lb6\�t�	Gz^R�t�(Vlm����2\j���G��1��
N�E�8���S�@�Pf���
���y�N��:8������= ��҉�?O�x�N��Ғ��9�-a�1s�XG��>t�ۗ��߽�diyiV8~M�D}�舖�+��!�U(��z��������?��NW��
�ǡ�<���_f�,G�L�#�_7�b��z�(��R$�T|�`=-�l7�p�,����{r�͂�,�<١{�<������ūX��~�����OS1c�4|��cfg�`��A�̝�>�>l�����?F�Q0z�a��Z����t��
�Q��Q��ߟ#~�Ͼ���k-���ׅ�]hj��4�;�:	/e(�J���)�L�?n��o?������մ���W�q���$K*y��)��@Y����)Ʊf�t��J�� ͎�Q_�\�z�?sā�4Ӧ��S]m?<�:^`�࿩��b�Yz��E_,��X��xH80�- ��?�Ahn�V�p~�QD�VY������3B�NCJWᥝ���F�giњ���<vQ����k@���6�����4=�O0Vi�fdI7�,������L�.�s�5��|��erx�9�vy�f��m�,!�Z�<{R.Y���׼,��,�� }7�$�~zި2�cZ4����'Bͼ�d�nFs{�0���ѯ�b�ٛQ�S�ax�>ٷ�ݞ�;�B�B��_qVj�;����ߕ`�_�v��k��]r�q@�������Λ�N�N���%�8��N�|�2��l&�h���m�dϣ\Z��S���� ���c 5	7��p����<�S���ն��Q����{��0S�Pk4��ZR��̶e����Md㯦�'~(�,��"}��"'8���Ȟo�8��H�8�H(V76��u�rn�I��<��8`��O���F2�Gw�3���1ߦ�5X�1�<���C0���m��(.��L�&�3��ޭ��@�<5��&��X"��j#��Eҷ0�����M��(�I�a- �LP+�$ƕ�{�ݬ-?�����;6tJzW������w<v�>7$�V�j]�S��9T]Ω���:A�:J����M�$�՚�mBD������ɮ�W��Z�p��SF��%#UJtV!X 	��c�^`�ML�o�B�NR���/��vV��r�2����n���O��OX����u�|�O�3���B�|�9m׸[r-��Y��$0��oc��|�S4�'6�7ݣ=���y�T�i��wF����O:c����0�G޳�)u7gX���v������&K��$�U�$�P,�|ث�z ^Ȳ�}c�ÛtS�|�Tv�*��gy��$���������/���s�5��"���߉H��PS�)$:p��j�3������D����]�8�լ����Ģى�pfc�⮌]}�5�dţ���zؖ!�~/��-"�^$�(d��o�'�P�7 '���}�&�� �{`3�e2O �X��'����]�j`�O�=�(�ʀe�������F���EA@J��{19) Ô.2�C�О�ޤ��=�E9��>�1�2���F�����B9g-�KP�6���,�CH���X���)u4�ܡÄDW�U��Y��G8�ȱ��?zj�,jtŚEғ 9.x3�Hm���ɘO<6<ٍA�&n���g��m�m�[�c�;/�bj��2)����i����-3���_UH�ӐG�E� &��G���l����mU!S^{nf'3��%^����pسo�)9�+��/�qٰet�V����Ҿ4@�J0��%s�E:8��I���u3���	*-����9�0��Ixt�����XOKO����h�;A�k��$*�"�b���V�/|��p�[�	���c l�EɥT+r�R�sh�|*���^��_�S��lJ���m�B�JS+i�#��� o���R|�^*����x\�Q����.뵉p����5�Y�n(�f��j��Vh־�_�}E
NDfX���3��Ŗc�O���3\c�c�}� �!����������ծ�R�Jm�A]�Lm�<�k������p:f����9B�O�7M�� ���YS�^\�v^�X/�j�ȏ}4�`�"W��4q�Sҽj���]f�{� ?D�1,��<`�G�����ƭp|��X¬�T!���ꂠ�r �ɔEjMBߠu��oT��j��br��F"��Y`���*�I�²��1x��@�X��]�#�R$꘻n�K����j;~�����Vo��F������E%Fޣ��-�NʆZ��-E��.��8��8B�;��5�f��e�|%ǂ0��Bߢ�^���d�2!q�d���bשK>��>Bv��V�!oŚc�~.buCNNOL\�����~#�I���h�52�Ք@0o�k��Xj�wU�|�Gd�N�k y�*c�UX*����OU1�f0��䳢ʂ����ф����o������N���{{�9a�sAC)�"Mts�4H�%��	>�6������\t�>Ͳ��G��܌��S(�~�0��q5c 0.t���G'��N�S����`�����k]�������;��o�x�o�ҁ��hH��l���ƒM�ۅ>��X7¥:'�aXp��IM���������8h���86���%�! �^�q�F��0�p�����eN�����ص��ԉT�5�Y4Тk�u��j�7������M`uݰ�$��ⴾK��4�j��<\�BK���aen��W���xм�W��Eȅ/��%�*Q
T�5����b���[�~$�.��q������|�l(wC2옍aIl��剓l�B�-2{d���4�n1���Vr�$��X	ѽ�wэ���mIɼd��ṍP�>r����KG,ĠM쐅�:�|����� �Oq�n���+�=tp��a�̨�a��6ED���L���r-+���H78�}�?k�g<�b�Q��#��~��log�L���1Ȁ9�������6	����5�%�*V7ݐ#�\m���Cn"�C��.��2���s���Y��XU_�j��@},q�' V�	�y������e��z̮��`xinUO�A&��w�n�5��!͑�7�VT>�G���6�M@@	{#{茧w��w"��Oo֍��K�잂7#(��xfq�V��~Bqu��該�W8Ѻ8\�8����.�*�lV����s��.��@�Sݑ��p�0��I�-ar���E���T:�v_φT�sT�ʿ]
�����V+z �y/S�����UvFɟ�Sa�}%T~��t��Ɍ32�ڻf��M��t��?h��,n
���B~q{�=/�>�YP�+��(�	�t,��:G�&��N��~�Wś�v�ե`�_gN�!���n�i�}�g��W��R���~�_Dj}k=RvW�X�_�!F7��բ���kKv��۳�7��/���^o������� թf�|qu�u��,k�+$�!�+w�2��[�� _G��t}Y�&��F��5���::�]t�>�@��d��"&����<Wﯺ���GV���IV�M�����C�U�v�xC ��l�*L�rǥ��̔-�!�ݥ�����>�#{�"�)'����):�KU��^2"���bL�cERH�n��vm{̔z$�^�R���wq�ش���B�n�#c{T2�� �}J2������)��c�c����g�n=K�B�r��X��4�w)F��F��'��"�N$SI3G�tY;~E��N<m�/���Z�!��A4x5�P�){�p<�{de�o�l�����:�gmk�����|��$�QNGs�+e9`>k9����֠n*��#J]�:C�9ft����vC��E�Xɉ�rZo�Ws\��'zX)���������1W)�J'�guS�~�(OE��s�<׈���Of�3"������ٙ��C�=E�*)s���,w\���/6؄Q��ܩ�������&|��	td��Mܥ���F��H�\�b�P8j�!�V��<��KE�6��P� 3(o��Z�͉Fqy��)�`��2|m��UtU�N�S��846���H�2��fɿ�d^�#Y��5�^-��%o�D� ��儚�$�|c�f��5;��eO{i��%�x&���D< ��5�A;�R��r�"ݖY^��/��K�i%:�����1d��_����gK�S�����h#C�$Fg���@R��s}r~�k���a%��6Ǝp��1��x��VЩV����,R9��J��y+�M9	��d�Q�<ҭ�	E��ٮ� �䏀Y}&�Vñ&3x�M�����W�Yg4���\D�=�}�h��z�G��b����j���da�X��}g�@�1�١Z��.(q����Bn'Q(�q�$�������&��J��W}O����^F�څ�Ki�6I�p�=��� ���)q�N�(��%.� ﻔa@c�r����'Ӈ^�-�~e
?Yq}L�Ig��K� ����s���Pet�΅�?�QkLE�$/QOpGt�`$i�[�k�����MR�z��bS����^
P�C�����Ҽ��������E.�[a
�qFd�Z=�yk�E�@������6n�K-�~��i��m�9��0�x2��T�٪s��Yb�6Lա�ސՉ�TI����Cn��g1c����O��DɷE���<:e��@T�s%I�I��&�?t���5��C|Cxb�)sg#�����D��U�"싾����=��I��ш�]�їH�����
n�`n9X��-�*�3��s���nr��1��9h��{Lj��0"Lf����_D�R� �m�w$;g 1ȣ/���j����Ke�K�+�����]��CD�u�y�.q��K�����-�������Q�г�4�6�'9�83*x�N6V0dt*0u�3|�"�(�?wX�¨���7��5������_q��5
!���J6(`���t�/�f�>�[6]/�z��M�O�f��=�+�Gmv���U��bޣ�q��g���;�Yo� �D	.2�Cx�aǞl�|I��A,9��~�� E��(��5¨��|������6��s��N�}����ׇ�hQ��D�O=n��W�OP>�A�� 9�uqB��g5���-�E���S���.\��[Ŵ<V��A\�3��ޯ�}9'��&H�Jn�a���H��m�����n��wY Ix~�.�́���	X�ax���rm?�u<�1�
D������	��ߣL	{�!�C?Ϗ�ݲ�Q�o�£CuMv����\���ٻ��{W���e��Њ�I�H������}ٽ�o��TZX3��z��d� �z�1��m�S>s�����U�UĲ;J%�2�\8m� �+$M�`:�9�v�DU�I�T_�,.�H�|���olI��I�N��S��cE�������c�����K�ZI��b�d�X{�<��p��=Sʸ�X3t�*��A9��~E�<�q0��#��T���T.hc[�\ÝS^H���b'��U}���q���(yY�>�%�B�>.�?���N�y��\�cj]��r��P�h��wǼ�	������}o�� l��s�T}1��L.�D��%��J���T΍ |v	m1%�aI�BAz��D��:�7��0���D�>�����G���[�Ml�X/h�>
+�,�����f��`�W����@�k�놘�����1\���D`PҬ��;��s���d��T�6!�;�V��R~΁��[�Y��z���cW���af]�����$^�sy���]w�**m�ᾠgEٲ��H��	�lY:�;7���y�L�!���3�j���Qٚ.��~����<:;�G�e4{�=wu�*\� �ՌÈ/�]su�������h��g|;���+G��n�@��j��b0?��~��.z�9�3������.3K&_VZDk���K����n���:��;���og�8�EF��3��NZQ���E�?���$6�>�9��1���/�G`qކN�	1�GB�v��e��0l/��ٿ��z'�o�(�TŞ��9BU3S�+�����QM��O� ��tk�Y�ov�1d)T�{�������E_X�$�8�,]�k6u��bBM��}꓄�#_�n�w��ˣ$�xe�N��Ћ%h�i�ҋ �8\&(�*#����by��ڄ����>�S��ܝ��Lz��ۯ[����y��Æʷſ��'�"��f@�P��,���d��=�q�=��B���+�UiC-���+4~�0M؛���\/tze�aY��畭���X��$���*fK x���̺��BI���*Q�E�9W��K�����^�V@�n3nT}�Q�a�� 6Vm�YH�fQ�@�{w�����U/b�(�y:�V/�`�*G7��3�91ИvQ��C˜��,�t�>h[`5����ך���j�sR�	�V�7���x�޲�r����
��*ox �[C��'�߸��3��J6�Ϭk�w�/I��o*p?���z���Y	vt��Q�|F���u��z.o��}oP����_X��-߂6	�N�����z���F:��� Ѩ��NZ�F��B��Ll�S;�2;]�T�9��{�����E���a`
o=������J�4ܩr�cw�ƺy�W�wk���cY�"���5t���f�f��%�r��q�1O0��\��lj�m,�j<�ҩ�ߺ�9NR@0��w�M��@]~ �_����������8�n{�M�h)[|bF�$��ʏ3���c��i�1D��A(�=���~T�����Y�4�`s�!����Id��.h�U���M�{��kr������%:���A̲jltϛ�b��;�3^�|;3;�-	��ӓ��e�,�Nr��g���q8r�&/�P�A*'D��(�	H	����q �yw���њ�qm�RfL4i^e-�/3�mg,�,����E�G�����m��5 /���t�獃7��+$+
�:���T��8�*Q��|���j�g]��&#��/M��S�x�����M!��/��uދї�u���BO��1��/���ۻ$ܤ�+�ڔ!�*���Bƫ�e�O���>��Dim��w\��rC�����WAv�\]��R� x��� e6��GoA��Q��{a��/!��R�e�s??�yё?@3,��Tt�x��gX�(w7���E���u~9�nI�^j����������t���	C�o�J���э��D�,��S/υ�8��]�t��x�r�Gk�;}��M̓,�X�ʦf�W ,��d�4PG%�Wjܬ|\ȁ�f-�����+���T��ڴ4�S��)�����ՊB�)�S���4����:��Kl�3��#*��P.'f���f�w(��R�f[���0h0t��A+S`�����N�s��y2z��{D�M�݁���2�1�dܴ��'�Buk
n/+/��Q�Q0b��*<�}J*Ȳ�k�R�\Z��/���	��		Z��cgk������S�-��Y��cp`kIF.��6�6 ���>�����)��*��r2���^l�
CE�-ќ�#�۵:��	᫘�Q"�A��F':���#h�������=ڿ1$����J�z��{�ꋦ���Եg��r�Q-|��qO<�1�SZR����*e���R�J�wlVn2��e{�¹3�A�x�QT��G��|("��I\j8-�t���[�	��,���8'\�U��qڡ�?���N�����
cg� �5�]�PF3sW��ՃH�[�������}�}*EWv��QP�K�ޙ��(��,��>�F����*��񴦩�ܢ9�3#�����(����[���3�����90=�,Nl�5��DZ�����qA(�\2�7Z�@�y��c�Z@'D/��	�DX�cЊ�y⯖
��m��P*�@;� J���"#s	.��ϼ�<�f�]Wh�i��l�BJ��~�k���Ү�+XJS��p�#{��CQ��vK�Ok�h�l�B�p�_:P6��ajw�����<U�����Q��)��3B�s�'O��ԅD���	4���oy��'H�5`�/� akG�8�:�FS�-m�[�মp|@N�K��*��m��[:��|Db:�j�"IZ�NQ�c�_��v �b��T�=; �6����=�I»��d\����K���
�x����vᥲ�
-�����0��+`�U�C\�Ͽ�-��I�N�X��>����@c�t�kTy�h��N�N.⁑=�ZrPuٮ7���2��N(>R�CbQ�/t���U%���/9r�����U�]t����߀-W<���}�k��~��Z��������sCm�=n�� _]$�|�����H�-#���ᯍ�ee�j7u|��\\
�S���~ձ,��ٻ^Y]dȧ���PϿ�q~\ �Y�A�ŧ����3�=R��'l|��V��O�h�-��5�ڝbT;G0e�;^�.��x�I���CU3̅�|�He2iޑ���������)�ڞ��~�X�y˃���.�8����e+b��M��r�����r�'ܴ��+^���^�����y���@T(`�y���7S�Ecw��!~2�+W�L���a!!Ԥ�U�{�7*z�',|^��]�����-����nEjo�RJ\���A�(�2R���tu@�s�C�I��ߏ��aI�ZK"�A^�w�LcFd���°q � )N����9ۉ�ޯŦ�̑�d6���f��|�U������
X��c�� �3��f*��������Y�{ח$Qҙ��}�zM���O�������7
OV�� �6}�?�^�dK�ٖ����+��?��:���kt���#
O	<⿼ɏ=u�O�g�)���i㨛H�D�ο��lऻ�T����� ��bM���((���RH��=Z/\��p�!�|����z��J���hh��o6A�VF4�A]�K��J'@L.Y%'l�r��o����cPi��6��QO�#�])'��ޖ�[��FX�;�|�ף&�v�b��p����cE�9�:�!9,�(Wt����i.O��sX�g��=�k��`HC��/Cp8��2�^�\�U B�|���I�k��j��R�,}¿5�/vI�]rD�
��N����ZRR؋8
�#8�@�I'��J1\ ��l5H�%-[���I�ßz`�Z���F�5��Lϡ�x;��r�A����%z����g�d9�Y`yH~x�����#�_dTTp�C� M��C�[h5|�f$Ơ;�T��O�,-���H�O6�د!W�~���Ð�7��J���oިp:���r���,5�YC��}����K��
�Fesb�qr��J���|.V�O,�v���;����"����X�'y�x��ƿ���e4|�O2|6��@��	�C#?�,՘�	���2[ڀq��j�B�BM�rgMv`h���E�>�Ҭ���6X����Z�uޗ�
5k���`[�o�uk�OI#�Z�싼c���S�J;t5�=�Hq��~7�~������7��T~��K�A��G�h���������@�)�x�0'�S��|�W��<��a��΢:�B6���r%.^!.剧f�i	U��E��K:7D?�~*�K�(x�2*��_����J��/[�Rߧh@�6K���`�}9����+M�ىK�ߪw0��$�2 :�>�]Z�#�%݊/R�qD3�7_zU$������r�V"�|S��.��̦:4�?j��s�Q�:>��������{ S�K^�=B�:z&]X��Ӫ�JiE�D{�7	yo�,���g�?u�
ڈO|�FGd�J{�h��,�T�P��Y5F+�.��ܴč)㎬H���:O�6$m��}:���>n������ePRk�����<��Sj�������g7�Gz�ɤ�1Q��n�D�pKRd��U���~x	tj�/*.]��mv�`o����#|v��h�+��XCt��f��)�rk��5�~2	ޢo�	{�T�Q8��!M�,35_R_�7���@)h��&��do�m��oRH�вo1��W�Qpgf������r�N侫�{�~�ت9"^�%d%�����GTL�qw�����,��{e��ݳ������!u"e���(��� N���fS;J�Jt��xmD�o"[|�7�Y�Ѕ`�~ >�
]zQ=��a;rv^�G�%]���u�����?���6�<�BD.ڛz��Q7�pX��� DG@��ֽ�&ܱ8���,s�5�����?�|�8T��-N�v������tܪ�0&p����:���¬��8߹��\�ă1&c��{��#OܼJV�I"M$ZtP/n����7hk:�V
��Q;W��DD�u|��k���L�#Ea��Bh�l��ڠy�P��l��7
�j
���G��@�'	�]*�%*�t���	��!E0�4b�;w�ǈ��τ*���(#~�`��G��2]=z:�*�k�.��h�
�1` ��Ԑ��w����L�)�T��H�m��%�Ë��!�^�Nl�6}p�x��8(q֝>BT�=ͼ�g>GuG�}e�쌴a�bꯎ8�N^"�xFiY��1Ju�oB�*Mc�8.+6�=����w�F	*
��;��d��v�j�Oâ{��K4�a8���N}��3�'�+��2��@��3Z���x3P)oM���@l��_��x��O	r�N�w'A\���Jڸ�d��O�Ј��jR�2Ƴğf��.Ԥ�΃U&�{kvG\Rd�D�[��SL7����k���˴�x��%l�)v�z���S�#���3�P��~�kN���>�#
h�!J"�;���8�odÛU?ff4�mU(��[�0X���F�0����P��O~��,�B��);�q���G~�?�jY�����~&����I���w���c�0��X#y�7�Ͷ<�� ����ܶ^�����p��^��:
������YV+����z{��M��������X	^��I�P�u,�i���MCo}ޯ�2X��v���d�s2�l$W�={�s%z,���<�_��,3q�'p�!���И_JbD����c#���d
<MΜ0T�)��.TK��'��!��1����Y�� qVvP0�� *���]���z�Ƣ�PCd��(��̡	Ȏ�ٰ��l�x��
�~���wF����YM2ʬ����q�*������u��g���[�� ��$��n�kfЊ�Ϳ��ʼ�M_F���Z����%G�pj~�r 05�����ä�Cn/(݁��Nl���˸rwZ$���X�a9KV�&�%ą��2UZ��(U���I��JD�c�����e��rҿد^���?5L�)L�vo{'�ߐ�'-Aw���?: .�io����e�e�)7�g�q�F��v�l I7�FV�~����F��"C�N]�Gɰ2�$�>�㔶�X�C��J)��2Y�9������J����-��~'���M��͂�[+��N��J��w�>���a��x�>r��ȹLo��5�˳b� P�T y3��@d����I#���6�M��f��Re�Ab�O�H�2D0��Z�1�����pRt�$�ҟ>�T;�vox�������}d��(Ct��d��-з��}�~v!X�g�z��܃Bm�ݹ�c��n��؊���u�A����K�)�٤��ю��[I�[�9cC5i���dԲ%̲���s�����m\���O8'/�i�8�)6E	�Ʌa��'�Ӕ3X���{���!}a�m���1
��������-��s�G	~"�>�v�A�u�����-"��B'c"������z0^�����BGn	�d	�7��ܷ�h�����&D�G,R��XG�|>�^Q����"z��Kf,Ԉ ��Ko��:���4���
��i|�OS��u�i6���4@9��_�\}e�GH"�)�;���5���� {~���EHX�:�M�m���3t)��a�c�nѾ��ʺ��-�:��dV�������슾s\4��$h���ae��Ρ�m����8-9�5{�U)�@qh���=u>�<�7mr5��ɮ��:�&���M?��&r%��fu�|ߢm����s�\b�qO���Rվ�~���D�c1����� _H?p_�)`L��h*��,��M����d���i�w>��%<��`+�kJKw��L��d���;Ԑ�>� ߑ;�wNr���b�C=�����f`��*��qa�8�v�K��	���b����@�4�������"�jK6e�ܐ/m>�w�6(c%=nK�кe�bAO9�A�'�$�u~6�(4�?B���dmv����*\��)xϹ�r�@k=�|N�3^\z�<N�)=ϛ���. ��.zE��;����P�Q6�F����xbr�n?$Ų��H�����R`F�O�����@B^��v�c�O#2� �4�ta@� [)85U�C���~�i�§��� BXj@��,{����`�QU�JQ�ư��ʆ���A����H1�;�`U�gS��ԙ�z|��LĹZ�ҧE�4�x���u�ܡ|�h?_�U�x�͆�F���o(���I(�7�[��s��]�Y�A�N,!���䷋/�y�˥�˰=
�iM3n��w��o������q��0���!�,>hAy�F�<oМ�2�!v�.��"4�x�:Pt$�
��di�?�c��b�@;z��?&�B�܆,	�f�<J����JV�<��zp��#�����Sz�#����t�6���K�vL�➤	��|������c������Z�椝bX����*�� ��"a�X��!v	���2�/��,XB��(�M�x|�_6��ڵ�p�3n�G���<3ם�Ʒx�����N%�r�"w�1�!r���'�+�A�|��܀z���Oyv��I%@��q��!.�yj�1Q�4�H�P����kb��Υx���$��-���.�������¨���J(+ƫ��Q@�ˣ����q�v k����_���UR:��Ǐ�;h�6�S��S��3Rl_���WM��,C?�oٚ�'�0��{wB��q���k� 5OOU/�Z@�rʟ_	7\��XjY3�������Y�
�k?'����a�`���0�2|cW�'� �7���Ę�CO��9X�x��H�[�\���b���\+�A61C�^���\NU���:������IG�r!Fg��UF���_2��������l�1��M��9R�Z�H��6Í�������yA&f}�;&d��d���"xx�tfp<\]��A(	���O��5�b��Jm��C��
�Gޏu/<�#%��'���KB��"l��@Q5�YF/"h��R�4IǞ=6�h-�
�k�V�$l��/�rۍ ���)tS���̡��E霌e���cn����d�f8�T��|uk��@x�pn�ҊfcRV}3�u���(^�E0A�R���!wr�!�#Hü"G�(5����t0m)+��0��NKЪ���A��d�o�չ\�ęw2kZ�v�
ΰ��D	��I�݂�H=s��1��&٧�n�C�7S:�Q/�o{�,B�c��\"Y�{{+�:����S]��2����4�������za� Y�Jۑ� 1�[<ѽ��6�i��F�4=K���S����~�Z����.��S�>!�r�(XG���A�D�-ۺT��	
Ⱦ6�
�����(�q� ې5dJg��i<=�J_�	�磪�r\�M$D�/y�.�w?T�.H�E�۪#c䎊:�4���n�ƴo��@�1e�G��\fD��B�\�����M�Aia][��<ib�v6�F�CdJg��os�2[�V�����`���O5/���Px�UIq�0�"V��概7�O��X��9C�"�V�Zr�J�U_���G�0����\���f4�82��3���]E��4E��o=���6u��*���<f��\�/������ѣ��`�Bt��-��V�U��ԩU�S�!�&$t	a���j��8[��v;�>����26�i�b���:d��aϊ��b��"D�{s�3�o]{i��j�[�n;|�y�]$v�N\��яM�}��|Q�p��j���1tǎ����J{�d�<F(���E����@뀦Q�ڕ��.�����6�cS�#ٲ-2俽�k�FH�$c�3s�]��7m�"�{�mM�G��w�T�p�����4N�L�섅{��7���9�>/���n,�7d*l��5d���to��*���6d^��M�?����X$�>�,��ëW	hC��M,m4	�u����1�kf�O��,� p��F�X*&��Z�x؛�h*���$${lϷ�?�)'��#�ː1�g�T�JX�&�VM���5/l�Jx�e���U���g䚔|/��-R��1�V���};}�HV���[�yH\)�	�,P3C�/F�_m��ϕ�Bg�v�@w�ߔ*��M��kq㫕���ĉ�=/��]��֣�T,B-̡#׮\,G/ ��E�ќ��[�W"z��5�|�{,���k����9���CcY���O���2s��_�`(�C�[l鼔1��>�<z�L�����k�m�|y��\#���e?\�wj�65�TE[t�E�y�6�)0�'�?'륶W��x-ow�x����U(JW����+��*=�{�P9f���k-�Ky�IJQ𗹝UlQml������Qե�@Z�J�<�E@VGV��'c����i-j�J�`5�@��Cn	a�{/y��#r�*(.��5�4�RE����|`�?�JA��f~�4�0A�����#�ޒ�,��՞��+4�R6�f�" ���f�A�<Ca�V���f-���v^�+V���tEaߞl�2\
���%*Y�'�x0��?���=%|dx����x��$�zj���Xl��g�qč�Fp�yԢ��>�q[��Yg#R�;e�C��+l�;j1�Bg��o��rg�Ӆ�OW�1�I�Vm �q���3!�z��!R@�⻲bzv���(5�E<ߍ�MT���P}ȓi�>s�*��fd@�V,'ʕ7�;�������je�G�+
<��F��E�@Y��
����Z�
���~�x��K+�˕��[AGS��˦Aao����N��
m2x��ֱTb�B�A���A�گ��GC\G�e�0�}�s�#�˪{��	?A4��o��}��
��x�U#p���h�lǂ���kv�2�XcL1��"wFat�s���AJ,[�L��0ȟ���Y/���L���v���O��OHS���I�$KZ�0*����f�������*��9�0*$�:�Z���A�,�vB�P����K�u^k���������.$'�H4
���p$�X�P�;�K,Ŋ'�[�B����߫�5���a�V�^��t6"�R����t�v��)o�%^POwV0��|;g:�p���i�>�g2Pon�/y��PbX�	\�9 D�L�w@���1��Z�\xk����A���Ҵ�?��АŢ���J�B%�T��q���E0��k*y�`.&��Ѧ�-*��j�o}�i]���;:�1Z_]<8ce3y��xp��jT���0:��owߒ7�%:lv��ɅNA;"�JW�vg��z�L�gE@=��w�����o-����F|6X$l>U�x:�u��7Z�\�OȢ��i�	HĆѭ ��{�o��wr�\J���d�Ԗ��TyI4{��W��>�~a�� �,�ixnRB|_��Z�S�H�և�\�y�~�j�&iH���'���RW8X9K�7��nx���xa6�I�ze��/Av�A� =g�����6F�UJ/�k>��Mfna?�:(d��?a��
]-�1�h�� ��`jn-8���K��˵Zu0u����c#�Qg�+����Or�a��w���;���>����~\��	+`�ݯ�g-\4�h�F���-[�v��c�=6t`Z�T������ȳ3�&f���s�p r��.�!2I pk�_fŬș�̖�%�Y�.5��T��ׄmC�����k�߰��ˀi���_��LY��0oLԻy^@��!�Y��Q�	YnV�2��zq�m��b��;�N�Gk�3�q�|�2V�Ŋ�Ȏ���$���wu���Pg�;�sBu+/]����&YD0�d ��܆]p�E���&C��q�Yt$�	#�c�2��92��e��Fs��R� wcH.��:�I���QF�3�"7�'���T9ݵ�)A�ϳ]�E����JP7Z���5�/���M�-]� <�6�q.�I}1��Y�����Q�[�`i׬`}���S@�9I�G|�[C��Z��0�Uu������K�1�4^�?��1!�f_�j@��u���N��T���x#փ�g@ �G����Հ�81�,{P�RlR�ıN��C;E)J�6�Z��Iq�ݧ��Aوz�gP��$�s����6��hW��w�����>i��=��W���)7��RO��#��	��LӤ��s8��RN(�R�����U�\2���� ���*b��=#����,��&�Dy�����{+�C��|��j$6��'>8K	G����p3�vn�'ێ�k�'��W�j8b�m0pɹ�C�8���ɼGՙV��5y[E85І�ESz�g'�aA_�_P���c��o�-���-��{㘏�*�f����h�r�����R�1��Tf{�K�2s��#=,�m��8BJ7�;}����4�l�)��N��~ Ag�tn@b��R�y�F��&�a�X@5}�*_V�q�E��A�>b���͢��]��o;Z��9�(�����Y��A�7^	���R��>�Þ꯹��� ˗bLJ���^�c�6n�r�d���cJΡ���p��ac���@�ȹY����j,�ңP(��K&�[�>���Ɏ����&/�vhx{	h�m�vB5�E^ �d�:(�tܴ��^+��%J3�Pp� ��U���e�������O-��Z�a��XJ�i�rc!�v����� ���w�J��*�n��{T�s�/v�� �7����q�y�4$Wn�=������+��j?yz���G��i�w���5�K�e_��8Ђ���k�}<�yme��fX�6���f<�
���&HR�C�I���V�5ϲ�E�������,߸V&3��7�2�ړ�Z��v_nL>�OA��s]�ʧ�ŷY��&�Zr ,�L:�p%Y���|�:���z��M@�P�y<��]� �A�2��D�+���3�bu��
w(��9F2|^d�4���C�Fz;�bQwZ|�uHjE�Hŧ����Pu[����5�2�4�Cj�|"��Q��R�ϵ5-yl�?k���t<�&����Z¡�;GU�Y��o�'��iU\D1*݂,�B'�yS�	q�WR/N�R�N���2�VgG @��P50�f?�F
\c��Z�ty]���zЈ�4+4I�3�Ŏ��2�"X�-i'FB4�����:���Ζ0�U��i~�w�}6)�����Z�4��;Y��Uzu�8�m�,Ȯ��W���,�u�ع���������	k�
��IGVO��˷+�$.K�oc�X�p��9_��6s���ȅ����Q/�~ç�'c�˲:�#zY������4|Tu~_��cp�R��+����2(�n�+�0�T�|�հ31�����7T\�~]���)�&��FgU�]�cQI��X�qk����8�{!���>p�Bj�nw���{IE��"'���&*v�d>3��WK����Y��5��R2f��^pf�/���P=�9�Tx�A��)R�9�yw�v�R��ؙ��.jÈ��Q��s��TlCa�N%n����!�!�����'���4���砂V���Zyk�����CǱ�}��K4�1��Z:�+�we:�9Л��w�܆�$��0��( Q������P �"�RV˵ggc��wnn=��R�	[�+2y!�Y��ygxF��G&?��A��
}�z&"�'�l0sM���1�n��#��9����V�(�rGx������d#}���*Ἦ�%@o`��wBݵYy���E�3��h<܆���4�XF!w`*|G���ᐩJ�C0������-̜�DqD8�{������.s��K��C܍MA}���w�=3�>��\�����~EK�T.���f�r�Q��C�;���r�a���Q/����FW��*1�~�,1_�^@25fˈ��O������Ef��2:��c�TG�N���6����ܖ/x�����+M�F �#���М0�r�\@�͸��lh(i-�|����']�V�I�r�(����x��#�uؕ~d��ZR \׎�r�PO������a��mSL~үb(w>���yą���v�2��wb����v�Qe�M�\�r>��z��h9kw�o����
����0CfT�U�2��@i~f�Q�]��1�%A�vN 2;�E�Twy�a���G+�N\؏\	�JB�%vJ9���?� ���(*�J)�Xt��c �.�dk�w�>��J�����@�����j z��+��2�AU�\��J��p����Z'	0B�5�L�
�m͓��@����bC�� F̗�Fs���j������HH	���l7�>�0sK@�.P����;�GB�����9M��o���G�����
��4C�
v*�!f��&�Ζ���:܋;�**��p�d�GЃ�\^��>,#x�Fev�����QC���R�!���B5�l�}�����j����X�`?���{��L�x���NR��´c��F��1X��i���ɱQ���VM�`̏_���B�B�ò�F$��#��x�I��,}�ΜX�x��I�"�����R<T�Q�*[��AQ6�>��L�=kK*�{�Hf�es��: ���`~��V�hW%�r!�ہ�4w*��w`����)1x�'M�_�a/z���
==
��>%�U��Ya�/�6�9]W2P��"�ۛ�������dOP�jX��߳s�T���r� �)q�}
p����G��y����%B���a;��E��5����iKLE��p�U�Z]v��m[�h�P�����R�H��:E~NW�v�6��V��Va�fN��c�L�9n�)ܑ���4��,<y1"�$�~�Y���Q_Dj�����U�������Ոa���́~Z���a��dz��A��~��ʗt�p�Q�-�D��
���o;e��/5��X�X��s��C<gltP�N�8�M�o�(DBZ���x�r(�!ʀ�UO�.��m!�@[�%H��p��N�h}c@��9d:B�˗�pz��#�&���̅��!����VYh����)ϒ}���V�!,�� �V�H�`hUS`_)n4��$i��y�KhJG?G{��(Se��$��!�y���2�m�������ay��Ƅ��߹i��wy�Q���^�!)�7�W��|�o��.�_�#8�����j{����n�y��'��_	��@z,����G�֧�X.��~�zI&%�ſD��+�ӊ�Z��6�����:��p9�]I���G ��v���-���sz���/c1�:Y�q
臒�m��=����=��zS����E|Z[hO�=k�a�
�.?�-}#�k��K�f�����LgfjWSЅ)���Xe���J�� ���eEc����_�Jm��9�!d����"�%��A�iべ?��E�bM���5�9=���%�VK���7!���p=�B����{�h>r 6��fU3UR��i��Լ�5s�'�'d=�q�zPN[μ�l��(B�̓-�Rl��N�Tf��W��I�vŔS��B�Po��E�-�a��zđ��_dw�r����a�e� 
��D���dj��k���>����5�S��zk/�f���.��t?%�x������ȓe�w�=�A�U���ی�;�ݴK�T扅F���k���5�'�C�����=9�'��Cڎ���W��Wڌ$�����1���ϡ��:J* P���<�V2|-+}�py<22I�*�Ģ�n;��Lbx�S>Ƈ���;�d�.���L@�����	:���0S�G�j�4zK�:�����aˋ������1�	���U�u�v+3mbfc�"҇y[�f�K�a������B	���kY�Y�$b,������OÒݓd��+**��D��@�S�R�o �﷼WZ �*�5���sx߂Ip�y����4�B-�xg�߇t�{J�ci!G������>��j��(��N�qU�g�}�A&$<���;�S�[I0i�C��Kx���R��@ܝ���uvq�q~D�.s��+]QQ��{�E��9�Fx������dz���P���=��lb�#�@2S[���l���r�>�E����5��Mz��԰f�d/&��4%���N䎌
f���Ü��|���
~~�a�rb�\��QEӷ;����A�T��Yo6�805�|���qr��%Dh
� �Y^��u�im�.��Cޮh���1]�_}�;R+.��/�j�uG6b�46�%lSgФA��s��b�d���9�V)E����iQ�eT�ڵ�Φ�Oy����@���0b���wQ����q__�~��FA\F(p2H%��4hmڄ@��U�Re
G>����<n����ER����,Wh�/S�`�V�m�-�$��5�ـ�}��[Y==���Ҭ�,���Z�Q0�6a����q��/�̌�>���SK ��k)�ݪ/�M���ܧ������(�["=��S�ڨ"���X���ҙ�^h��p,��}��m���`��^4E�Tz�~S��OY�Q��"���Y(-���Χ��	x�6��A3�F|w���,�`����q�w�������8��ص).�%G �ب��Ib��h��}G4��6��B���b�I�1_5V_^�n�[ŧ�����V%����!�M�T���-�'����T��tLo���*�-�f���ɵ%ai�U�$"kkr� e��*OeA��a0�a,e�h��/T�;���C����Z,��v&�B��f��^��[�Y!��k�+��t�-�f�a/����ipDy[Z�2yR$�V�L�u��L��������0N�]g���#�K�Z�$	9.,�v�3ɮU/׫��Έ�x�q�I��(�'T�MG5���)-������e2���}Z�� "�����^��q�2).�.B�i� �� �m�4c�Anl	"l�LN�Z��0�v�ޑ-���������{���v�Z�C�_wGb*�U\�}��qQ�S)L �ٴ���d�=}�׋n��.V|-7tފ<��[�ȝ� �ib3S�0�.ö�bB�4�ķw�n!�t@��-�[��]���ȐI|Y}�hy�Ĥ��ذΉK��iFC�7!4�/���+�c�g�V�1\�"F�q"��C��wζ��/�-@�6u8%�|<z�RqMo���3^G��J�RG�w	�U��z-yt��$�u�[ ���=�H|���s[�|b^��;}$k�uA=�c2���sI�ԋ�(`�5����h�}���A.6⨘0�n�M��撕q��|&�Z��Rc {t?+!Evǿ�h���?������/��2��v�|�ƩV�H�a�0�q^�+�X+�XO�{F�Ǘ�%��:�m��B ��.�]xٲ!��)Y��R���X$k�c�8� �WKG��3�����t�%�
��\��K�o���]��Lh�2`I�.|�8oK��f�v;��-Ū�͝�K8C���� �[Ŕ�ת�m��O��(K'�򙌣�Q��~���¹��

�h���pSk \1[��תn�R&af�R{�*�@��\r��	�/��;��,l�S� /h��E�s8#N/��{�C��=Q)��f��k�I u�pg��2+�9T��+�5Gj�¶)�$�h&�o�)�9�[D��T'����#b�?���v�DI��w̳RN}�_8�%�]u���'�m>K7 ��S����(͖���z&%�-�x9 ��d\�p Y��#̹���@TcD���L��,�ay+�v��:�`��Bw��H��-�Ղ4�BAѸ����r|\6�H�fzvv�6���!71�ܡ�����W_��5�F���(.�~�m��(�"��#*+�S��.PZ�����m��ӻ����c�F��M�đ�sV�J�����P�6#Wa[������Y�̠qZEF]�{4�^��d��I��l���2H.���o�����>�$D_-v�����������m�x�{|3�C����mN���jKE~�Ҥ/�)��L�c�	6X?��M|�����0���O�Rκmk�A��VdC���r(�- C��fTjr5j������-؁GA�5P����
��@T��2W�l��:�� r�t�Au@��������r}b�'#�,�&+��j�3X��	� �����W�l�m��G�=ޢ�NB�HBA�t��_K%���a�S�G��Z�}G�����b��諁��[9܄�ߦDN��u[:��s5E�֜�H�k[�Α���~Q1� ͙,�;,���͌��W��&��$�H�7�d�+N�3��(f0!c(�N9fV��&~��1m�q/|�/5��SS�7�����|����g�Js���*��3�K�ROtr�$�q���8�-��|�r���x����h9D|s�3NrXĴ�ՁU^#�@�O7���#/�\�.Zp[��|*o�rS�_��F_=|!��7
|<W6�U^=�O$G�����! �U+�ƭ�̥l��&I��'7��^@�T3}ݺIy0��;�C���9���	�N��5 $��q�����c�B__/h����\[r��I���,L���u��eҐ���>��q�I��!�m��ϑ�;c�ȵ)b�sݜ�@G��^� :�<c��6�I��gV�4[m|~x��S����u�E���3�-o����\`��Z�܁��ۛ5C7n6~ଙH�ף�P�� (B8=2��fo�"tiB�,�<%�j�8i;D
�
E"��ۤU�s�
VP&�By�ɫ� ��sn���qG�gk,��x��j;�k�^�b�k��Dp��l:J#j�X	���9�v��c =���[5�;�i�m�"��(#,�\���L5��)y� ���	�-ui�p�2
&�����Y���%K.w��'�y�: �_Q)MG�fkn7���;�t���yw��r��D*Ci��T���}��凌����;߶�iZ�,m���"�!'�"���7���m�vC:v�h���"^O?�Q�g�!�j"��hEA�+��K�e�Z�R��^V(��gZ���0�BYA�E!6Ο�>��T��#�{8��a4�:�ɼS�4�����e'��RG�V<�0���g�,�y��/�B�JhzH�q���hL8@�D�&��M��䜨sVPfx\\�mRN&�)atm�,���Q�����r��`�i�}%��Ukƾ�}p�#� ���l\�f�Ծ�x���SZ�=_�]ߺTa���R2�������K@K�?��Ց��S��Tw�^k;���[�uX��FV���y.C�
��ZOehu'�O�ƈ���vԱ�v���ZԞ�~�(䥡"9��h�U�C~E���D�/+ot.��XZ��NP4�dx�Hߺ>���^� ��9:U둣\��n|$�`z��,�t���zخ���"��g&?�Ž17E�X��<҃��*/|90=iI��x2�w9��/Z��g�4�L��	A:fƙ����Y%��[�33)�/��6ۃ��:��j���)cTv��hTq�Mk9 f�Ϩ`�����F?��쒎M)�2;�
�o���tԻ,n$҂���=�PɒLLO��EEQ>��Z�6����e�:�-%%��(�U��l���A�����&����ț�I�T̹���ΑZ1NM]YB����Y� ����V��C1��B�hr8uy����(C��)�+��+zy��T	�P0���`N����p��}�2��3�SO4��)�m#�)f�K14N6���ȡ	��Q8����ht����c_�QjK14Sn�p��M'Z��Y���H�?�$d
	ix݇B%J��~lֵ�p��`Bw��1�$�����,m�Fo~��!��$�i�S78��)+w�{z��w�[�#u�R��ю�W������WY��ћ��e��9A�?�Ε�y�E$	�`�6�R߶3�\�cF=�u�gI��o��������N�Ie���Qt��+ٵ#��Vӕ*s�"{��]���`'��X���S�&~�z��.�ɜ�T*O��?�����B�^�wZ��XIM�{���X�I�)r+E��]��#9�4���p︊�aM�E��T.����[����j���V������ԍ�:�U���q�r��<�m$�8O*�������xf��Z�		��2�	g��wS[޷�,5��%���`�]��k��1V��J����a�]��mD74
l5���ǩ@Uvn�X}B�tꧬK;���;�qoH�q�}W_1�7���Ia�-����70�`�㡩�z6a�ۖƮZIcn�k����n<�7�� d���gkJ�{�h�n�cͱ۠����l趤�=-9n1Ny��w���U��z+�����J�J�TkG��AG zh�>��N��kO����w�y�=�b���"����[�Ԕ�=�����n�y�=�t� BD�C=6���"�jF��֝4��F|~@�>�g�*}|ǲ
�c�,xE�@���=q���P%λ��`Z�7˔�. �A��"J_��.UU|�+�T5�����q��S��$L�7��]���-�yU�z9����ƏVd�8�l��a�ʷ���%I��Z���{zyu��#8o�]����{���E�ۚ�e+�._`?1���y�w4&���j0A��Y�J�������sؠ����,�8��V;�8��d�P�u�K��X�"}p�g����׵0�,{��u�QyJ��3\��aX�*��������Ǫi�#��W��U� G<-�1�+H��򨝉����`Bդ���9B�Or�>��c��̻f�uF�p�%+:��7�M��I��O%�����-�8�g�
�ъl�����k�<��/��`�Еxk�n`i�����Dn�\��UWŁ�	��d���g+��#��a��Ʈ_�#~M��ev�إ[�rTwn�)�]>��-J x�[��NWb����d����u����X2u�mGr��=?(��&�q���.wHP���������p�R��N�[S�n����-�S����T[�a�yXʆU ����I��:M[)�h�>/)g�7~:��z�͕����P��}t�/[F�-�����`�t?�'�s��0E�N�H)����(SRsDK�S)&�Ŏw���MiĄ��Sʌ�O�Lw�4�n9G՗��p��V�Z^3�����:K�ܖZ�$_����y��5329iXY��TE#P�l����s�b����;����6J�kj`,�|��l�1�p���,oi6�PH�-�F���rs$��"� X�?w�G�y��_���w���L��r�B6�j���Lt{;i�������`�Zej�_��H��^�4u�q���GF��U�*����xY6� ��?��l�{�"��`N����}>����|��	�^��dl�&*��Q�A� ���CY�Fmr�W!ްk�Ձ��;���[T��~�+²ك`̳v*p�"4�vԺU�a��ڙ�f���O�`���I�
�TG��̴U�yV��Pd��"�~|�3�� ~�F��Hˡ��3/Y�#��C^��j0#<R|��Dp����L��~�־+]/)�p�b/�l��G���҄���c���}c%:f��J;�	(I�#@&�1�x)D��� ��3�ݏj�{D��a �����J�[��� ���sv[����a�z{�DP�M��Ô�L�~)���G��GBA#���)F�"� ���'x���g�U �ß\*&MX4�M!D@���{��S��(jv��IL�-z�y�d����@��@-*�20�`V+��Y�	9p�$��3A���p�j�ǋ����뙕�H�V'��?7��TC0�"Y��U�T��<�n�A�Fù���7����� w�,��@���?�ՙ�ׁ����Lt�}��?A޺����a���T�� 
va]ILo�cŪ��$7)÷����� �<�z������j�hǬp�j������u��m/�n+��H��pg=�GKy�����P+�'�kP�j��'N���f�Q���?��o�qyPץ�f��%9���R&���Mh�Fd#p�yY�u=^3�Nf�:3#Q��u�;3K"�U
,s����U:�0,�'R�	�/s�
z��2.�}s2��q.�T��@��I�Wy�T�uc�1`X���E9$��' ����\[��Y7��&�O�a�~*N�+���hb_���5|�����|^/�Sg�O:\$o*��>� A-�]ZX]0Q�����SvV��響L�����#E��i@�?D�7R7�(�|����z�}y�ӨD��	ވ�[y�|��0#�<��r|�!���e����*��[�Nqvg1�	�cZ19����/g�n`?A�B�zB�ل?^B*�>���f�j=�4$��yӟ㲙����ֆ�Y9ǚ��������4'��0�VbA*�2WNV
��7��_Q\�6�)�o�#H��]㉲��`?��!)�܆q�D+�e����T]iEZG?ƅ��@�qy��-���<2��T����B>�rg��_ �������Nmw$�.K	Q�
oI_��_��U���[J���*�mQ��s�V������N3Py��3X��A@-*Ǟ¼�6�<�8�N�<:Pq��S�u1�|R,K�B&���FhM���^�G�Y�o��6�*!sC*�G~�k֨�Q<�"���r�ECv w[����k~?��sa��\��:��ݞ �S�X���hU��a�r�p.��8�ю�E��њ2@M���D���c�9ıS��,P�l<�=xb���ӂ�PB�Se�h�x*Ѵ�ws#�z;�Լ��骶ѼPMOF1�����[+R�$��e�������T�BI��$Ip;4��M1Iz�U^7SY��.��*����-5~O��=�0�1 ����ʮ�EE�@ņ��,�\һL�E��>b����J]��d$�IPz>�4�ND�*&qĊ�_��Q�dD���!J� d�Y�ĜV���D�lїU�Z'���]d
p'�aM9��w���?��h������^�VƬ����e!aV�z�33�V�t�-v�yQ��������mL;V��S�RDO��y�*�aH�<b�m��8�p�`>R���w�l"�V;��V�]d�ʫu��()̭�\O�$T��G-ogeNӮ�ݥ-��R���m̂���y���q3�=��c�j���M�36ʉT��Fd��	��]n�q"���g��ic���R6-�W���>Y�����3-�~�H|�~��e�/a:��_�!1ո�:����@����],�p�|I	�r� u[�!	W��n�U�E��q�<_�n+��")��ߞow�IX%RB:�ѷBp���2��p3�F���f�ݕ�E�?Si�ѽl�}�%gশ~j��ؖ��7����`���d�v�?�"@�R�������o~��u=��
~�ceJ��s���a<���K$m^����_��h?���N�X��*H,y:<��d�\����9�]�*C�F�r6����
�')�l�aҰCsd��hU�*)	i��T��cv��),0Ed���t�p�V/v��Ƭ`fd�k��mh�^9��}�u�o*�l5�t��S#�+홡�PLy���jL��I��0���)�0�(/��0Z��$v��]��i����K�h�P��>�����K���t98[�ƒa*U���`x�����S4ǆ��H��ig�$�LE������3�-a^�@�oS)�g��Fi!���]ɢ鍊{ϽU,D�%��rYKMՆ��&�0���=CO#��MO?��޲Z��lȲ����A��1��#,��@�2�1
Kh}yϬj1z{>����Ք���/�6�u�:M*�(���z�k��N�l׌���W��ZT�ų@q�T��L���DPy�a�����w�=����5~A8*��A��������*��dX�ǟ����%*�0g�']���sa����|�]j�>  ��1D��EI	C�DdzU�A��+���ٻ�:Q��Y�yk�?Q?3g����\�Ѿ�DR�K���q$���?|)�Nc�� �MX�+j�yD�_?�?8�� Ӳ�%�$N^Q���j�@Wůu�3�ʄ��hU�∴� �N&���Y0D Md
�MG˵���l�Z�4���������T��~����?�v�zP��ưQa �/�r lBx"�R�i�{���X����J2�(T��Y�
�G<��5ټh�
�������9�T���&ע?
�_c�Ō�8��U�����B,��S����d�,��S(�V����ӊ��d4�z�u��Rw���@T��O�����-�.�~֩ͷKq޻��]�Ib� ��ٳ�٨���<�#�^�OVĶ�8���F|�+"H!���G9�b(a��b4�o��[�kv�M�D�K&4���{5|'�@�y�����{?��zL�%~����3Sa�v�*RLb"�Df��Ļ��Ιu�Q��Ѽ�C�oB��V�Ӭ�`�Έ�e�W��	(�軟3\���:k�`D�i��N��3�+`��[�'�|�nv��U�2P��k�<cF��� �����o�W�>5���?�h��B �E���n�=�
B@5�82��-���C�ⶖm܇�b�(��p�+��tw'�}q(�Y�W]uD�E�5y����������z�� 8Cͧ)�vK����r`��
+{�#�ܝ�������d�A�
N�0#)"��PO���:���w5��L�w�S�&�	�	K+�T��!�z����¿�&�To��ϴ >��p��Rp-����y/�cAvË�5����7��Qo�}U�]ɱܒ��r�7\X������l�?L8-�)y�G3N'ZcR$���*O����1� $��^���t~FiPU���ܛ�PT�9�+�,	�[�<q|�?^X��}n*i�����[�ڥ|ơT���~ٔ�]�쳛�o�,�A҈U�S���hz�v�L�0(hy%;�.h/�q݃}	Q55[�<��+jk�t��M�
f���A+Ix�u����wK����z�?u��*E�T���ǌFG����E�xr"j��#������3ͧ��&��&��!U�)���[��wS��e�ʞ�U��yaF���ԃ��*N�g�����r9�y6r�W��lb�Q3���?�k�+#|�Vǒۋ�+�s�̟O%��Q�{N; ]�î?\`ղ=���H)J%L��~Y�o�L��E�����:p$ZU<�]�������Ȭ �&:�Y���o�Y�n?���;4����KV���N'��#{@��3Ey��KNU��T���V&� 5�a,)��AV��f�ʲ}f5�b���#�o��BT�8�D�Uu�6���)/=�8�*m�d.�
~5(��kԌ�O��ւ9r��@r0ڣY�,��v��@_�͝L��e&4bt�A�Ǳ�8�v~���A�M�iD����]�}'��;sY�H�e���Cϥ�|z>	�'�62���'!{��[S["z�q�0v,f�ך���ϟWJ����ex�1yG�@[�����*�8iD�����.( ��Rhڲ�.�H	|V^?�X=U�,[��Ǯ
W	��s�JBT�S�.�!>�����_�����?f9,���pӲ[>�^�,���u]�bĵ��*jTʵn��m���;K��e8Y�)DL�c��ݯwٞG4QwV��}0v�"�i��v�S44X��n�y��\"C~MB�X <+"��i-�x@Ǡn�;�<��r5�fU�5.6ˌ_� n�7�`u�
��;^8�n�1��㷽;8�2��E���g��Tni�H�[��,��ݸ�˻�' ���?�q^3����ҤeE�����,H��}��>�gM�\N�P��O0�����c�ٝfv���~�du����@ �|��+��P�!ʽ62���#h�T}��U�ht�����0�yK}52m��jKũ�"uҞ` �y;���� V��{Y}$�qQ-[5B� �h�Rr���yd�tV��͙�~(��,�c_�D���~��VG�����o��:yA���/�'_�s�-e����L�w,v�\`G��/n��NU��"Qq�k�F�O��TB�~#WwB��a��b{���E��[���)K$}T9���MSg۬h�N�I�������/ם�0a/C��PaO�����[���&t[ۏ�뺶|�9�{��9w��z�A��"�,�������:-L�P�u�|��4!1�+�yJaB��-�>�l$�K�QYS�1	�h҆����T��ـ0F�^��㇯��%�ᘕN�W_>3nI��Î�^�d�����pXm6��0^�#{�w��uca�N����I�����h6���2�l,$T�4[jw���TY�@�q�,�������?�7���x	�Ajfp�Ǡ�q�_#�)�QZ �"�?2�A��6ܚ/���`\h8t��4�Y��{�_����.�m�S�y"�>�K޲j����ρ.�;x����}�k@��S[��Rqh�l;q�\|'�~M�c��-�[sUf_�������N������u��?V��|9�b]B�$Y:�A-6�sc�`�)����~�U57��-r�3'<�N��/eJu|�!�c/�WNA�t9�������r���5"�O	d�`����%����m��9�y{��z5�f���1J������\�<��2�Ձ�(C�{���ʄ���@��2�6 D������Y}E��e^4;�a��_3�|\
Ӵ��ۺP�1�� ���<@�rJy�g�~��
^�������P���#}= Y
!.|� r����t�#F���*�����D.��7/����'�㌗��2�.W�.?��a�B�OM�6�R�L�����g��!�r9�p#��'�!�_@���r�{M��K���	��^*z���3��皉�V�~�r����;�ga`��-�%���'�U������,TR��A}�a�	kEt�5k �W��D��W�Mae#j��|p'��� S�6�����9����tu�ÿvgS�Sfxhq��| ���u.7���_�$�����P��w޽Ϻ���Ϭ�Ώ�h%�u6�CTs���T�P�@�^9��YhL>�.tq4�$�|������1�*~��}���K�3e�^bgy�ID���(��G/���ݡ��4Y�Y�[��ݤt������A�捳�ר{������R�Ǣ�o����$J�8�:� ���j+����m��Z�{q��^ȟ��k���z�����^��01����|#�V��i�k0�D�fI#�<K��j��C4���H�H
��������-3�8>Xh�����s���]����P̶*&�-��g;>a3���O��gURtZ�¸I���<�x&' ����6�V۳i�d�Bd:���ӄUL���h�Iw���=��]c�?a.fe��6�ɇe�C��է<�3w1�����K\�C"v������p�Q'4�	JO�t�=E��rl��'`z���߀���3sx:q�t�t�c%����ʖ�=��L�B�E���s9h>��j>e�E������U�W�YIe 
$t���C�D�P]]~D��Ĉ��L�����tNp2�y���F�`Ov����d�y�S�p�ɦ�.�d����y�,U(�}�C��b�������b���%��cM��=J���n ]�Q|��N[���A��Hb�ћ�
	�n�|m��K����1kȇ-ɨ��Ms���X�!	��>v?��M�x�(H�J<���iU6:���?�yS����5�c�Ϊ��_���V���6���ֆlN��J�����Ԝ)p�ha��0;D�c:�5��
?�<�-�v��_�FN�a\[9 B��y�������SBƚ-ޗ��"Bp��њ��P�#4	�	�o[�I6ny@���CY�7�=Bz���GB4�ᯥ�?��X0�g[`g��������rC։p��7��jb¦P ��t%�[�A�1?=CQs��+{	t�������]K��ɲ���g�Ӷq�,Q��UXh��Q|�{J���s���v��Jt������\��t��5֝�U�n�$�+5n�H,���N�Aԟ�������� Ԡt�\D�@�k9�U
�8=��;j�"m�w�������>sdSx�S��GIu#0��a�HV �F��+��3���q9�������VS)�=����S�h���ܗ%��tr�nPSsб��*F�pҠpE��|��]
m<h��K!9�����.�����Z?�3P^�6[.?��1��M"��.���N����̯����8�#!�}�i%�j�x� �' ��-�5�(<��Wׇm\��V���k#��&��ϓR��.���������|��,w-�	E|��`PZr >P�
���ܘx�WL�>�P��U��&q˂�έ� ���ʸ2��Z���bv�l�6��_}�OR������9m��B�u�n�@�?Mhv�����8���&]5�4��}9ѿ�Ƞ��D����c�O0o؏I�,��{�X��@�^�Pc��w��::���EI�Ή�D!J�ɴ��%�j��S��l�G���a�t(����r�s�V�mG�R9�F�m�i�jtl�i\Z�����)�D+a���h�E`����3�rqث�T�WPwM���h�d��4p�:���� ։�H��0��N�Gą~���o����{�� ��6@n�9_��E�kǦ�̗���׬4���g���粤YD�I��t� L=#��ryԥ7:g r$��:��w}<�j����ՠ�%0K�ۜ��r�.��>��Gb�}x�Z�=�)s���s��&��j��,X���J�����,����`M/�0R�l��#�Z	:;���2M�+-p��?	��V�O�
�r^�S9�keQ�S�l�G�=��]Ü�*�N�/�rxm�'��~U�r��������X�1a���{��a�F�<k���LQ�Lq `��fw�k�' -d�㩎E_�W&�.��>���� ��JQ��x?'[+� �y�-]ǯ�r�x,G�Jm,�z���4-X���x��&D,,�p���d8ymD��0��q�[mΙr%CsHp����f	Ou� ���+�����>[��B��.]L�ө_b�Iz�����o�	��~n�Tk�.Ţhh9��Z�^qX�v$��l��Њ �L���p��~a�Q�v�D�7��éC���G���s�8���o���� 8f���V������%��7��ɫ)��glWT�֮��������\Aδht�	`�OQ���se�q�
J��6	sk��SU�QKRȂ&�&ӾR��K�ȞEu�I˴r����^����E��n�[Lu����ќ^�P�L8�<�+0�t���=h�z��>6*��K�-r�v]�O����ۈ���'���1ij����3����̽
�I���k�'F��
m��ۄ�<u���S�d"���m4DiB�ŝ��tSg]�׍�V��:{��V�F�?W4Y{'�t[��� t�Ph�=�8��Qk�=�6�{�JY����.��螦�6�a|�Wd�2�h����t�#,�X�5.cd-TT{���������\b�fzT��7%�E�@mI��y�����]�����>�J?r&(*f?<��H-Ǉ�L�V�V��QY�Y!��QD=��ƫ/B[�����5�WDr��3߅��(�2&�־{�(|��\_?ܟ��ED��]{�p�x=|�C�����!�
�q̲�P���?X�{eJ?n���+�^�3R�6���7iw|�
�;?nnP]�C��^"�9�gs깱����Qbs��J��P�Р��д�	��Kz!\�Zݥ_4{��l�OWM;#g�=xN�:�G�y !�d��KDRK"u� ��E55��G̕Ʉ��}�NT�� ͭ�rbK/�
��#t�x��b�#�8�`����3*_����P]���\y�iM�~m�k����4e��+�QQ$��^e�h+L>�q�Z�b�g��GT�s��:�礜��$Mī�M�=�	u|PJ���:��1��G���������բ�oh���j��2��C�������$DG�nJ���?�[��_]�*����7��ɻ"��� :��e��Ov0�]l��<*�!�w��~�?�[9�f��M�VsQք$��:�<��ֿ�2*_rJ����ܞ%c%���X�o�K�M ��'��ٺ����pM�3�hp�r"��?q��.��;~�����[!���{���� �jc"�E��=�L�fhسSebE�8�x��k��g�L<U�ޙ��3�}�׺}��F�����g?[c\�x ՠRଅ`����� U�$&��d�26���Q��p��ws�.
������	���~_oI:�!$s'�"�ɺ��)��6I�T��Ɓ��u��z"���c��*�$D t?5�5ų��Z�kj�9g��*�D�1^�k'I%B����D�_�;TR�Z�.l'nvc�f�~�����#-��[)Ƕ+6��zL�uj���cM�Ъ8�g��pT� ��dK�����Ìi��?	�b��1!|}L�ai��T�;�h}ۡ�]xY��n���F�ֈ��s�����@���@9'��=��?� �>�>P�dl�e�p,������1���گ���.�|{��H,&\h��8>.�Z�_�⻳��x��La4	6U����/�H���5�����,��s8�\�Ӎ�o��uG�S� Q��Jԏ!XЭ��Yp�Y,��܏�l���<7���v�C�C�ޱ"���#Y�/ȃ#-C�w.l#P*��$�����_���PY��Iw�q{n���`8*�tV'IJ�����'Wrr8o��-G�@��9�Pd�,�O�Noq�Nabin��ܛ���|
��".܁Ώ�����XA�u䱘�gw��˝�O�9���*�6G�z���\��5Mw>	4��l���,�i�>�/�0|q~ss8��@�ܕ�uɪ�II�m�"��w�|z�ku��,���M�w�Q\�yOU�������t!��۠ds"�e���oS}�Ф���R�BV�ԺC]�+�d�BCQT��|������'�N���L'�����Ux�/��Q�y�x��G�Ô��/t�hZ<vׅ����4W�{ �]7��T��/Ԟ��mx��W΁_n�tW�u�M]=D>��l�6��o��@f�����椷�|�'H�:�ݙ����Q:��u*�W.�%�����2I��:YhP�+����X�YqF^�����e �Ow�_���j���;"�2
׻�������Q��:��Ɵ�mbtO�N1��sc���9P��f�>�oCi_c���i��py�=��M�)��]��$���&]��:�����C	K�~�4�%�@���v�m����� ����a0��Y#�c/������ K �CC��M�l :��cs��	���:#ۆ����������[#�{7)\�}�0�}Ȼ�ڟ���	��HyN�§�|"v�L�H�����A�t^��D�9�<����r������np�'sr1Y#)A���G������\ql�:�#������ī�_���S���kzωg��e�ɜ����㠈�%-{� ��E�E��gku��[� z��0�x�0;���@���\2�!��cS 滀W�nA;��h���^٩>ѓ�d���!��?���v�B�Mr��k��٫�$d��a�{>셣�����H�l��>E&"9)��rޱ�莠��Wφ��4K^	̱a%7FO��ϫ?���B�+,�c䌹�=���L�v�<	�a�����ӫ��a�@�B{�����ڇg�ƈۍn4�l}QU��[�O�T�R��p�ʘr�����^h�m  ��&��3� Y�#��/�{��M 3��������3�%�f�z����㜹^�D��#������폕���n��b�R�mvQ���5�%!�!�rO��!�oy�lh�Z�[�q�r�0�GY��z@>}���}�.-�?�H�i@��Žjk���@�-C���!8/M�Pe�=紐�x���UN4��������tC�He�U(�_K�bC���EQg�.ˎ0�H��65RVM�;�KF�^E�t2�Y���(�rC��7 �f�ֿth�>����q�M�E�����	%)7l����_G�L��^���!�w���_����Zyuǥ4�,;w� ���sR��%6�ٴɐ��,ʒ1���`���qV	v�M��R7�Ϟ��r�x-��ʷ�|[���OK.���>���#���@�;Im�������Ϧ��bv��Nk�"�R-!I�5W��&ɴT���>%!�\x�K���*�F�o{I��0���Ng=6��^�!~��-�0���d��e2W�l��1����׋�4Y���9w���۷�u{�7���3��i]U�3d�U����Uo�p�,��8.�<C��7n<8-�3�6��gAS:�6�d�����u�ݘ��t��Se���*W*D����[r	��v�@^��~��>��N-4E�|�1��:3ұ�#h����6ӊ��v���S
]��K���[Љ9�y��C�-�n)@�������vX�<�?�[ҋ�8aR��3:v��c��&�q9�9Ǒ�آK;*(j�_���g�GP�.�&
�)�F��DEla �(���0��hl�5g㤦�:Q���>7O�߹�.0ef~$3N�c�j|��r6�ܦ���E���6qp7�u:"ѵ0�{���%�_�����%6mϕ�g�ʔ�>��$M;���ɴ�����1�c�R���O��_O����8�� +�&��u�`:�v�:�K����NI�����]WٖE��`}S�F��X���a���Gm��,����hߜ��䊱[R����/��V{74C���������J���6z;�*ө�A�%m���ۋ*ّ�<bop`�1�?t����#BR�\�M�Z��h�D
UN��4]�hϾ,���"��Hq��D�#��'�s{����b��m��c�y&���(���3�M v��W}\�E��μ��Ϲ$���6�]�n�W%^.t���D&�I��u����(���g�\��(�B݌@�w(L
0�7�rvp����C�?FBw��E��E	�g!
��W��$d����yQ���J�Fq#L݄}H=)x�Ps�0�k�uTiaS�on�[V[N�?I�iF�C���agS� �]��4�մ�S$�{z�L�k�B͎q���d=�C]q�?�c8K^�ǐ��3���
r��J�u�|�h[F���P^u����Ւ���$HK1lu�7"W�I{�h����#��+ɏc�"�N���N
>d��&��2?%w��|Aw��wMRͥ^'XK��_�Bj����_0�#�`�a�ʃAR�Wm��N�����B�e*!�구߅ZL-��[���ν�T-]L&��m\��)Ga�g �����ν�H���E� б����h�a�	�s�C��d�<��)5�JG\�uNc@V�R[��뒉,uL����N�#3[�TA|[	�����H15��u��x%ᥧMcJ��y�
��I$N.C')�y�|D�8(�{�t��Ll ��UNl�������XnV�a��+�%\�>G�z`���t�D�t��i�t�\\G.���,���[��+ɱ��*�����+< �oJۃ�)�������kyH�ʹ&UZn��cj�Ԗ�˶dtJJr�jr�?/�5~�������=	�s�}8#�RU��|�L���qc���Z�m�ٓ�U��c���Vܾ�$xn?�y��Z��)�b/��:	�����fKˣ蓉�����OCZ`}�}�vsl�4�XB��P9�Nu�N��>2���:�FT$���6�ѹ���W��� �������Q5dkٙv'|xNÍ�����
>�+Bp��@P��h�h�FD��tgP����T�8s�C��:#�nv�[�kj8�EhOՏ��;����5@����l�����4/�zi-���z���7i��AW�O/�9����IvC�C����=^Eǽ�s e(JR
�X�g���@3�i9���\|�| �	\�[���i]�<z��lQcHӰ���ys���\5%6�v��g*���؜h�Z�����L2:Pf����3uI�1W2#�T6�ȾL��J����8*��9`�O�+ܾJ��C5q�h�rɺ�O�c�|�B�lJD��P*�a�H�=��M�Ҿ_�wP5J"��5	�A"C� ׈�R���M�F��&�FA	��[
i �h�%�k]�ت�:�WA�������N�40�/�*]�Y�O�Zq�x>�P�,�nE.�_G����I� �?�۬��w���ﯖ`j�𸂽E��Q�?��50?����u��X�<�F�o1>Ӟ{���Bӎ�p��M�d���^1Ŷ5��k��������xe~�>G��w�}~���r{ ��n�P��ũ�J��'����˓Ʀ�K�@*�0ܓ��B������y�ځ�$��|�����a�������x�9Yr��=��p.���`���']r��;���,�w2� �&�����Y�X���+���.=�Q��7����7����ӣ�<�Z�q�Y:���ՒOW&ӊBrKg;����F�76��rǗW�%���\���WK
8*��v2��1d��G�y�����Y����o
�uE���|�)1EO��A"1��O�M:g�\��J�@� ��2J��؅����)T�_�9[ێ�5�ʝUJQ���bH���4�#���[D��
C��)�,��P�o�k{��y�y�p��k��/��G��5CZo��f�7N��nwҖwD�O0��|�L���W�"�Y(��Qڲ&?r�D4NۦUj%�	 ��}Q#�%_��]��*u~�3�#X����C��N6�qmM����@�]����՜��o 5�Rh�y�P�dF�m��ތ �-=X3��WO�pUx�-�1G6���R��3�"�>2�Khz7��<�R��3�Y!�%ŴK�����������
��J�8���9f�b|K�a�&�q���U�y��e������k�;�afX�j�yó�] �(UA8�~��^����3>���A��`���$�p_��~�Ā7�x;'5I��џ��|���X��O @$m�t%OR���C�-�IN����g��y�Rth�����%�H!9=�䜒G C0��)��x�`x��Z��WG�ui�L��Its��'���z&��]<��aW��bQ���}0�)x�g`��u/<���fZUQ�p�L4���!��
<fV��heM!�F�qj��*U%B�3.=���/���M�*̉�>�8�����^����Z�2xR����ίN�~V&Y$мL���}�`䞌��JT��eM�|~��� K:z9<.*&���]7ی笛�¯�j���1@b=Ke��ߛ'��EI� �����=�|A�H�K�n��H�D(AR�=,z�o�������3h��,��8�ђӠ@���x���b�Ƶb�{j����BF��_lՅ
j|C1z rJ�����\���VlXf��ZX	��[W>�նM�5|�)�Z5z|Y&�<���iaR�4� ��e�4V<��Y���Q�3")	���A��J�V�$���S��D��Ì��|%�(#:z�n�g��yB�U��o �LG������_`0���Z���qQ�/r��i���\J��.��o�
­+_��Vah�OL��B�"�woj�Y�vK>w����<y�u������A.���M>�VojVkS�Wځ<�f��ǥ� ��*r:�$��,�F��Ý��?�qqX=-�lC�nZ��h�F �B[�x��h��HY��߯��f	%����o\Ԥt(��PF��h�s���TW��q��8Tu�:p��Pm�u�eO��$n)�Ib����W�%-�y����g����A����{E�;q��<9io(U+Ӧ�!/���B�d#W!]�<Y;�o�$�[(�<�O�<p��i��r�q��	S� ���-ʊ�o�E?)�ft�xF��jlN�4����S.#�|��űy/�#^�a����0�v�.�W�L��B$6��K"5�އ�O��CV�5/đ�Ay�=�V�~��r��z�ic򉼳_���@���%]��
�I�� �f�K�{�����;2ϋS�y�Ig|# }U;~=o�$%���qi&
\�l�Z�������s�8��χR���S�@gN�N�7� ��ylF��/��䚂�ɈG��uw�ܝ��.1��v���6�y����+��p����}ڬRKG<��T��S�ӐRN�Lvi.X�o������X�W$��F7k˨eH������0~�1��x�<��yrIg%���)��q�v��8Ƿ֒�f}�٬)"����=�}��$Iէ��U�^�u�W������
3HO��j�#���1�TX�A�]�����X⇻d<�׃���:�sM7�)���^��#�J[��	���Q gQ��j�[k�:�x���]l��v�Y�wSqˣ_f���t�i(!��.���o��P����,���l�/���M��"D�B�|����&A�������1i�^�7'"���oR@��s+�0��[Mr��5GW�\�&!���<d��N~5{�\S�47�����܋�F�\3&;?k��!��@*YF<�?����Զ��_��V��D�ui#�= VI��Z�<�G%Zdj�h���|a����fڊ�~. �(:?���cI�����W��U|���6,_*�p����onj�zҽ�h�s�+�C_�l2;�K�feu��\G�L�۰w7d���f-��Pb�Y$"�q��q^gU{�t�*$��ؐG���Y��	�fe��"s�]_�^�Ϥ�N08��KW抁gC�����Ǩ������5����U��� �+�8sF����������p�P6�r�iN� �\"K�n�B%��[�
V6sƔ�&�y�F�)3w� �pri�����hg��G�w��$z�'3FZ��&#�wL#7d��xX�Yr3��
C �ی�8�
6�=�ө䨬��V���@�øcM�okN�:{��i���3hV���4F�G<pߕ������!�OR����g��F7����P��е�[��!��[���^�9s�'���O�Z��+�Ó�8�����Яʅm<(Y�=��!2��v�z��+�=�`L[�?�aL@�b��b��(�*Ls�@PZI�Z�	���c���Fz!������"GN�V�&u�=w���Sধ��"0	v�00C�����4yM\���l}��y}o��6a#�r�.Jw�g�w� ��<ֳ�˰�;�q#�9Uy�gj�ó���ۡc�[�D/�ш�����Z�sO3�-Zk�P�'@Ɠ��$����C�6��2��(W̝�/�p�7���:#h�K��3��_	�F�6Bdޓ9�g���vLy�X6��2���2#��Ⱦ���$����]�$k]���{�o����y����
�'7�I�q�� 5hcM�z����4<�B#EY��֨M��y��;�!Is�����9�}��r��:W�>%�YY��,�-ki������~z�ң�|�x=���3Τc�-]�^�T��T�9�(+�:R,�"�]0��)��ӐetoZ�8����7�@"��8Лz �o^ķܾ��иp��`�M�=j`�ƙ����~?V:<�+�n��%s���3yG��<'�>O�ƿ`��5>4h��5�n�S�$T U7x%��>l�a�e�C^+NZ����ݗZ���Wc^�>�רy���}�x	ÞR���˿^bH�̺�e6S'����y�n��O�=��xF�r�odڭU���w��n�r���er��R͏����c%Z���L+������p[l���
=z(���E������ڥoT{+*H6�uǌ�o-l��* �v�I��0���	�U�"|� �P��R+4�eO��g�KQ�Y����4����x(�m��H��;p���gb�6zɳ�d5�X��f�gJք���0(p�,e/Ѐ��#����:5�oI#ѓ,�e��zf͚�!ø�H��JȬ��9�Oޣ��`mm���϶��an�a���G20���������!'�8���<����`p���]I!h0�3Qx����l�NP�l%B-M�rD�X�4��v",��#��$Iq~0]��~�?,�J��3<�7�a��D�r�Y���~��Y�L1`�il�B�*��"���W��2^�j����>���踡a��א}[%��>�A�`pq�f��j���2��W��t�X�.V;(>0i�I��ވek� ����U�x��J��S�q8m���C�T^����ՑO����g���lXT;��p!>汏f�dL���z�'��b7��Hg(X�+��W�4�E|�P�A�WNg�j���౎U���NnI���Zn[�F�[��J�t	��L:�qB���V�����s&Y���c&c���p5��1tvX_�;��������0>1�� ��|�3}a}V������1���{,�X����z�p_8�4l�/? �*���H����ݑ�,�]vbC)Zk��;����:��1O�`Au?�?le!�x{�{�}X7a��g$��)�1Gi��z
̀`�dA\�D�������Jxh� �Q9ѫ�"I�fs���%�G\ql�y�{d��V�A^��)��л�6��x�_|\���9)V}���x����\����͐y@~���bE�*=�g��5�ϺӞ�6�U`ɮEHZ�޲p�o�����A+˻)��X�@�L�G��B�!2^�k�U�l�X"���E��	ךE���E<uF-�M�l�T�t�N�,���'ԣfֈ�o�k���=[e �ɘǧeQ�P�t���7��'�u�������5=��K��H�nU�	l��H)M>�,��?�E����Y�<h(��65,WmACj��I������y�r��t����&��5[l_v?gʋ�	#]��x�v�A�	1�6�������vJ�;�*�R�9��
��.�?j�y�`���M��S6��BZ�o!�GF������R�d)�0�i��{��� 1��in}�e}<H�Mj�`j�g2���X��+K�+�h��M��j(!���~?���'��I��7d��>�qX =�"�T���f�i%����C��n�4U1��z�m[���(@d�C�_Fs�
0��r�]
u��1
�C@L���#�]�B1�ꑦr��Z�d>Q�|X����?�N�O�X�?L�������Ҳ	���508��h7�o1�k�7���㥌�rEӤv+�f�?���hw.�s����2��]H9TF[�
�dL�Wu��i�E�I{��(�{|�:�M�C���~���"[C���$��8

K�^/([~$*��遈��V�Q`���d�+S�E�\���4B��3G���D3j*�!����lz�ݬ������rߑ~C��M������0���O{�xv	�&ۂ��_V�#IcDb1�b!���l��=��B(�AD�Q(�j�X����u�25��v��y���G^�'=>�ho�~>y��q��Av,mBw�'#�ڲE^8�Ei��U{����K��o4�z���	��jS$7�9��0�y�C��,tԝ����O�C�4r
e��v(�n �\b��b�/��[���R�9A%��a�}���%�K�R�!�f4� w�S3���{xH{���;�۽�;n1��M!1��BS�i��>bw���?"��j$�!
������%�v��t�����G�K���+1ҽ_���v~����|#���L{�!��u��3���m�m���x�cj_,�{�����~���3�eu�[�Y�^�[��eC�X���@��mS����˭��d
�IVob=���!,�;T��X�d�O�j���b�ݱ�T��yN�C�$���r���K��7��%��4.��4/��� e�ZA����GD���۟�3k��X�Y�G��
}�^�+F�D��.k3��] �	��$n�M�/���(a+�<+2jl�ə�Q�7�x|�(�$֦��,��h:x�1~����)����E��:�t�Es�!�߷�N��	�����7���:'�]i.N<h��~�S��H���a�N�����E�p�/P���)�f0o����ݛ0�i�<���i��5��#"iv��[K��	�m;T4f1�sB�3�B�=��T��v-�"8�j���a������q�\��KN��>�L��aV�)��"O� րz�B-�-n��-I������z��7��Ų,�E�yTB7�PN�,�_�vQ6�[q��O�Ho�X&Ӭ���'!���Z�y8��D07�Q�߉��������g�M`}��?�e���T0̔a�y��޾5뚜�(x�Q�[�ٱ����TR�Dh�)�.�3Eķ<��v��~����2,�1�T�"��2$�H�v��uO��ʪ5;������eM��{v����h�oN5\�P�m��J�l�6��vi�!lÓ!%��n ��z�\:m+YrH$I�`��gJV�pa0�X�U�O TջE�Y֞a����<�=�5> ��G��4�|��+p�wZ.출�'�-2� U���
��ʅqǺ��e1���md!�:�5��9Y�+u��7��u����"O�O�dfM�H&�Y��zZ���W��lĚ����i&�[g(���(V��A���?uO��-���7����#�m��Ccۼ�D���OfD�6��RnN�$l�����=Z#cN5�x�5~�4x4R�耔�%��Õæ	��4(C	𮧑�x�u�&+�$�$��Љ�":����j��h�5cgW�N"��\��.��J��	3�.�#wm� [ʱ�D.vD
u��ԫ�i$ 9��|��<9�Z:Nkn�n��zd����h�Q�@�Jy����`�}��8�3
:�H�e�ht��UWh�}m��ǒ@�
X��q����?)�r����¹sۙb9r����.:���ؒ�AC_�&I�²��`��nX_�hS��6/���%�l���^�
j�"�XT��[�!Nq<��� U�a��>��D7A��S��2_=��z�_<��~���q\6n�_���p#1TI���x��qyu�1��@�
uk k��[8�5(�?�vC�|�r�/,��a������Q�[f���>:	d(8�#� �5��Y8N�h�[]�����Al�\����x��L�|wIw� �_�ŒH��l[`R٠�PT[��Ώ�(TѸ�w� �.v*�s���N���]�!�PO��m~y�����Q�!�ޟۓ������r�2w�:S��bL� ��4"�;������RjQ�£�h�V�۱̤	�ա��y-��p~�E
�G�m�9�e�;X���9oC~����S�T��@e�Y����ޭ�q�ߑ ϖ�+��T�kN���y��/�[�wmg�R�$!{<�?��p��5��z�=b]m��[�-_��C�]�\�C�ad9a�"_^d��PJ��ЎVdR����k��G�1���%��꜀4���t}�Bu<9,l5��>�@�i���:���z�G��4�����Hm�!h��-N� SA�E�n8�se�"R����![��=w�I�d%,�O~b��H%�:�o�<�s�WND��	�K��<�`�/������^�ݴ�SN������=��Y]O���&m��m WߟpN[�*U�#�.�^�����x���h�����c&:�i���ʥ��h�N������ѿ�6���P��,��Q�Xu���"�S�8�d��	?:���3��Bap�!��B]_p��w��L�X�]�z���i�V�8�G*�ߚؿs�ݞ���[�2��|����b,np�SV�v�a��"ue�Mp������=�+������RdJ6��t�e�0/�X�Ɉ/�M������+'8og�U�~Ju�.e�M�ya��?�̫�G|h!F}���p.�� ɬ�٣jBnJ�����.pI�7IIo���o ���S�Q�L�W�K	�� ��K���Ҧ�C�I٧�\"�VfsR��\vW��Vgn�׼,�4� L>�AR�!�3�_q�6��cR�D�y���N�$�����r3��5�t'�FZ���S�w*��"��J��Z�ez�mXMNcC��IG~��g7f"V�����
|�o�S1��`��~��ww ���ɨN���k�[��0o_�����g�a����w�ɲ&
����-���;��>mab�V("��Mo<5A�hơ�Ǫ�J³���Ag����}MV�"P�-B��Z���ظҒ5�G�+8�ż��y����S�	�59Ay�̯������00�j<͎@����w2a0��O}��B��]��������ۻ�|\�o�����r���P������Ȧ��{`����q=XY���Uf�Tȯ��Cb=D42e�g=�q�ASe��%m�z#�!Ǌ�[_�<x��i]��שv�	0>y��Z�M�l�dӜ�^]$�J���#ٖR�װσ�m�����l"�`�xrT��MEY��ȼؾ�A�i��8><��^�=`ƒ��e��o�S�d�'f(��r�G��o�S���%�E0e����t�Bp�u1?��Ǻ��oY]�i Q�D�����Y����h��i_4�7jh��
U��O`w=�I�� ۈ���r6V��-dV8�P�C)��n?�[b�0F-N-�#J�v��=U���տnQ=��la�z�m��3�����d�e*�	�G���t��TEa�����1)���磗 g�Z#jG?u�U
�u���"�������eg�UK�����G8��M� {3��Iڐ�P����f���%�g\�  ��6�.�	|����:�d���Y��'�c@y$|7���Ii���x���L�L�ײ$��V~�w:��:q�(5�w�jov�"Y7{AY�w�����W:3�H[�`{�
����"�vgw�Ppq�Z^МV����\Ї��ƮL��t�ς��l��Ϙqo0���
��O勰]N���z&�%�,/M�7�m��GRJ2�
�ҘLP��������酹n��g>���5��	���q������|ld���m~J�;١�<�#�[�2R�m�g�{��{��z�*�Y.��,h�3D1������"�QmOy���Q�.VJsl�Ѷ�:��T3�:�&�^F%_��s�����z<��&Z�;`5W#�]7	�V~���K?G�^Efg�j/��pX�]:�v���b�5^���#hV'�ZU���IQ��#����8wf�p�=��e�<!�`D��QS3q\���t����y��̍d�Y+��q3S����;�頡t;>	g� L�W_-�@��aV�r9�XYƗ�
�I^~��b`�
I_<�����KO[��
j]l���8���xk�_�'�x7�5��|�Bz��������#Q�lǆxK,�����MN��'����x��n��?$f�����K�i��m��+3�m>cC2K��)�!�D�8'��2�Cl�� � �����Hg����x����b��Qj�-�~/P��:_u�琯��*N}�w=ƍI��(*�ͳ�l�<�=G���[A�ސjBf�gQ���l~Z����C��r� a��40�J���g4|\ES�J��&�0�	���=j���岋O�r+1Ή���-�e��S�m�@4����H%Ą f�Iퟻ�g���* �D�b:�>����1��ه�$����S�aR��a$v��B�J++ig�@'#F��5�N� |�xCr���!��$͎���ks��>ݫ|�����w��Z�����??dZ�j_}qIv�<X`�<�yY��Tϡ����Y��J,��1�3+YKU�c����9��2���.^た#o�%��48ӽ{���%B�h�������b���Tm�F�|v�z�V`��hB���W�H�V�I92l~���&;���I*[p,�@�]���o �*�����]=jG���&���5���F�2F�2�]�+���0���!m�8��F�y!�؃��	gdfι���}�-kBl뷸O�(��Vp�)�+\	c7J���	������1TT������f'q�0�o�s�_ME����\��t��&H=�!U;��t���t«%e�0	Ɏl:ջ:�VC�aѮ�U����AW&�q� ���+X���*l'��?-��;͐���WT�I3\�}F���u�=^�q`���K��kNдm������O�
"�ɬ�]
�_�^eN�PE�WmG����1V���䙍m�w����e�J�r��c?k�L��� s��ة�u�\����H���v��ao�V���Ȧ���F�q�#M�h�1��󭘊4���=xqp:~���jϞx�e�%аm��#�'��`x? �]�S�j�|��.:*�^���4J�G�LZ�����r�^Ze�35sѡ�+UǞX�_�,���%������~�'D����/���m�˼�Ca�Ǘp���� l��"�lp�/e�e�)�79���3�s�q�6wCEnK0&N�}�Ղ|ؽ�<n�T�%Nd�.��r���'C�6��ӡN�n��]V�iZ�b��� ~W_��$�*}iE*�d=T��&���������w�c���lc���Z�D�qDt��Z�q��W_J�17��FK��q@L6���� � ,����zg�} C��`�	�&����;"h��8^�p����s���r��������,�h���4{Gl��s:�ϟ�X[�L�T�z`��,*�b�@N�M���b��&�d#5�)F�ތA!��?��+�ߟtDE���(X���my�k�������S]�I�(/ơ�}T�V����=�ݒ�J�aE�ܒz�<�|"�B}ܼr�7����l���/�����T3̅�N��ܺJ�S�XY0��/%�n���P�Y�
�1�_#��ٴ�{�FU���0�;Ha��&�:�����]���E���T�5�sƳ�)9�A�֢v���(99 3��џ��7@��y�K���Ev�x��	��+!��݇�[��5+�݄��c�^��������'�Ed���������c�kcp��Q��g.�W���䛝�	�t�?mP��Z���!���y��x�>��#�{�N�Z/����"3���\~��s���Ư(W���s|'�x
wD�k��{�� ^Զ���/��s�ïz�����`�,"F��m�_9x��������\�+ؕõ�\Ӱ'sU��a>9{>N}��{:�z��������KԢ/�*v��U��o���)e&�f�vhZZ�T��p��)��`+Tc�8��S�;�w����8T5��/�Y,�4��J�b(�t�)0:��ϩ�$��K%:��P)�mb���[ jz��f^Lc�P�i?�G��B�li�Ӌ��I�r1;�I���-f�U�ȧ����E+ę�l�e���׎q`1~_cD��=6-<}h�wԜ=���k�P�V��Z��y�K	f:����2���Sj�؛�v(o�8�q�r�у�@`�_����1�s��Os}�@�VG�����Pv���o�)�
�^��L��%1�˰W
w���ݾB-��k5�C�͎�ε�M��ݜ!�'������_r��q� ]��q�m"����b,@lB#�I���Lw�	C���r]�z�7�s^�<���]�T���tX�@d\��R_��*�3j�)ݡ ��޳M�;�R����;B;�|��>�F940��oQ���R�]�??�H2"Uۖ8���:���I�N��^'�ha}O�z��}yO�h�F�
?Z���R��<Rv�G�4���S-�����	�|P�wC���Q�<"fW�UG$���(����R��G�Q���6}x�H򈣆��>���4e4�Ƈ���Z��3����͹!�sb�0[ ^�L���[c0�Cż��\����1���5�F~EAU.�h[�ey�~��\~�J6����:ή?�vK�:���I����w�ɻ���4�{\dL��NKX�2p���k��c�F�!�=D�j_3���D����-��*2F�S�F�~�%�X!Ue������୿&��0��hH���[��Jaî�N�+�J��IC}tY�p�y.��&�v��̾�Pk������6�;b��_+�o�{�[��U�qc��튤^�����J��i�W{as&'J�s�8���:b'��U�s'��}�jê,~oL���q�@����"w�<~�I�JA��5�⡹k����u	�L�+B�0��r@�#�j�k�^Z�J�x�^�[,�Pؐhd0�/G�f>��1��l3ƪ�ǉKcZ,Bt������r�L$.�;6�'���?��#h*��	#��Fq��3=����E��Fp��h��������e�hjK�HKEI�� �]�
D�P=�%!.3*92�r�[�q?�Is���U&he;��DҬF{OYH�Uo���)���ޝ��|H���3��Bi6�{3����5F���47M�:�4`=E����'+��� �W�=��L���M2Vel<�TVb�bnEa�F�ْ}<����Ƈ�GP���Ϊ�s=Qt�G�� �ʨ���#˵a�?��6T�ӹ���wR�X��p�0��RQ􍶃��`c�5D��B2ۭ�����!�T�p�A7
�>1��x�[�X���R�J�Fb`�< ��_����@\�n����#c�
��]���cr�[����_����x�AP��n'������^k55 ��Yv����_�/�M\�ܒ��9bN�����I$V���]F#�:*4�]�m��y��֩�|�Fkt�A���g���M!\Dj��A�)*�JS>�������8;h5>�ƽBh��3r����a�A@N4�����*�YG��zG���(�3��!bI��*I���m�D��<Ǭ�_8KR����^� �l�ѼXf_���2r;+G8d5}�pO�=h�ͤt#��e�_f�=zCxˡگż$��8��%���.IHȇ��R�5���l�2����p�t��n0�4!�w����J�����.�����Q����
�4͎�R���Y �U���d�O֠S�}J�Y� ^��9�憺��Ҿ�.���{��@�K꙽T1���^���o�(F�[�݇e�y?\�r(�������U����-9[�QH!w�[��F��*�Ǚ�oW��+!�f���=��͙�7�1���W�_��'zs��Ry����)~�("1����,5�R�y�����ўWQ1<Ny{��iP�x�х��e)�|��\%�E='b(�!U���#ٳT�z���|�9�&���$�w��#�ɭ��񦠺1��ѹMf���	����j;e��<�-��-����C	*(�8��/�Ȯ�Ȫ��'r�]d��WI��2������?����E�C�k���\΀���Ž:��)���Xx"�̿�X�q�U�AȀ��]J{���!�%%i��o�jhO��e/̀�P�7QEj�Ƣ���,0s޹��G�T��;��FB��]�ߕ[Y�uw��J���^'��}è�YD&�rc+̊�\fö�.��Vz�"���E��o��y?� _�w�i?��Ky]?AYe�h��Ha�o��Ե�3��>nH5q�߭�S>���(�$�`��#!'a��Y����-o#��/��C���SU\�P�]�p��>Ɓ/�Gk����ŰO��k~6��į�Me��I���#=�?�6����"|�a��$�%
ov��қ��s5�C\S�B���-+r���_V+3ġ^3�R���׷��.<��<	i�@�d�^���Y_:ݏ���� ����+�����j�QV���GݢB�_<a)�k�p%<iJ�xg�'���Yf�蓎M�1Cʹ$�.��م}uj��>��N��2��lc�w�?��.#{��Q�N&b}@HX_��x��� =���;��0|mP��4�����^$��Ev�i/w�I?8��m�j������'p�9�ۂ��V�Z/ߝ������IuJF��q[a|��)����c[I�K$�v2ݍd��8����Ha��2ãq7�^�\��0+�|U� ҧA%�f�'�PU�ĬC����!8/����]�ᑊ��R"b�3�����{��Cb�+�]�0���L�4���yS�fY����d֨�C�"l��P��+�n>ʲ��q�=!�v�Li���ؔL���e�TK�������feR�#0��������j��?߅|]����Ku�Q�J� X��B6��Z���f�~2�`�>���A�}��<J?A��q0��%�ZQK$6�д�a`���M�c��FĵAs/��{�l�h&*d�� �����}�ܓ�A�Kt��p:]��=���m_��>�R�f�����<V��oB��P���`������NaN�v�i�K��)3��Ę����lk����>��e�$�狉r��.�×��_�����F����ޏ�\����;%_\t!��ژ���L�T^E�X�j�at�D�l�2�O)ۺ3W���	&s�+H^C�6��~�<����t��	@��qA�.خ�8H��Ŧ\'��,lJ>$�EU��=r�;��gwҠ?�Ի8��n��t��T9�dY�Ԗ�I�R`�M9�]԰����4���)���0��� g����pA�b1?P7.s5a�דpH�<QXO�,0ʴ뎷�fi�s�y��5�`��1���򑁃�C����2�@��~)�����{��0V���i�=�FO��(,�]B�� �\Q�0��{�̇�8��0<� �h�؈�<�����0fK�(8/��J��
t���Ȭ��6 �|CO��f4�?�涂C���Ñh�#CP-�F����w� aD�T�wxjJ�f#*`�BƢ���;߾��,UK3�0Je7[2�T{. <TZ��<'�8���if,�:���������r=�b�������6�[l����Cz�nu���v��sZ'f��+�T�) f9�Cٖ+�3/}{�R]�:�߾��F�=��ƛ�nZ��@:�;憆r>��Ho����oV���w�o�1C;�<L\��Cϟ/?q^�h֭���B��K�GwRJ��u�\Q/,�I��z�����Y�f�!T��)Յ�S=���G?��`�ֵ#�:̻�M��T��)^���.��B�5����,	�E�x��}��|o��J�!RY3_4K���Қ&r����?P��QiP���^Ppy��焬?MP�2�5��M�l^yW��_�����|dH ��PT�#�<gFis(�x�ې�(�<� �yyV�z��a�Cs`�BZU�� �hy}DP*��'���b�����=��H��댒l������7���!O#_�֟�0���Њ^[��`����ɂ$��1���[	����V���7R�Q��8VƆ1���3��-[,O�˖�˩O��	k8�������ș�I�Ka��A{��Ȍ��y����w (�+�E,�tX��e]�B�)��ȭ��>�o���
��YZ)f����F|�oME�C6Hh�}�[���%�/a��9b�'��_�<����Ԃ��G�71ږ=�ݽ��{��ؖY���=emn �bщf$�g�V�i��0��Z}�ǃ�7�P���{c��R�v�u�'���x.�<�y�q	�p�$���TJ����xSr�B@_��$�N#?��?-j��%�t�%�^Ү!>�s>��(�����VO�-�NE�n�V4qE���HͶ�e��we�B>q���H�!��v�Qe�u�"s'�w�V�du�����,]�e%���U�# ��s�"��%-�>�Ȩ�TlP��j�1�(?�V&��%(l�.�ڈs'�b�+�1%q�����쏲hF=�6
��yO*�UoD %�A՗�sJ�U�e�N�(1jO�#��[���!!0�R$�e�*\K\`�z�Oݪ�<��8
�o���t��ۭ�J�'�0����eg�vƻ)��e��O�J��o�+�Q���Rf+��*s4З5�)E�`���^�Vf���g®'�zZ~C6wg=x�/�YW�T� d�������B u��Ry����q�yK�!�8j@��=��b�����d�M����jc�#9�^|Gz3�)\�C)xkR�|�^��PIL�S���*��&�f��q'�w
��ح`X��8,��hN�!U�B�o"ɕ;�P90sZ_��Y��H?M`���iB�!-x�k����O��Ѥd��4��H��5�rPxq3�Z\lq�6����ټ	��Qo���L	�4�e�{0r�Pj�i�q�q��Ђ��-�G
�V��a��j�7'��i�ů�ok0yW,GI�����x�h.{�:*����2d�q�@C�L�M �|�+҈y-����'�$׫��q��%��>��� ϭF�Ԧ�J�'�Q�S�i��x���+����hb�/��Z.������7���������V�\�k���Y�c�Q�Zz��0z�F!^!��m���?�w8:�uCO�c��u��%O��.�g�G/'v�OC�b�SV{94w�d.��P�pP�T�){������Z,1�G�"
C�<���韊�YGx��h؀tE�窖}�B%k��"��x���Ѽx�EL*�3�`i�r����j[
e��i~��_u�wi?���'%6z:�7K7�#wޒ�T������p$A��q�V��2Ff��y��dK#�.zf�õ8��uM��l��e�r^�^F�?���m![��}��x͍�"�F-��R
N����+�rȯ�������ͽP0�w��f��6a&j�s_F�"y�T�:����a���[������i/�.q`g���f�or��az�@�
S_����ϱBM9�Q+{�<��*ZOBқ��7���fc���"ڤd)*�[14<�{ԍzt��3�Jql3�����yM����A|)p}�I�+>�aa�Q�+�H@�n
P����_(�(���p�x�(��ne���|'�y&:��d4�嬤���f�gU���캠(��l��U����)dup2=��e�9e����\^&�2"�\�4�PRΪ(<ef̦�W F?�$����Hu�BF�7v���j�T?�_ UE��{A�&;�і������L���i����U[�<˾�&c,*V;�{��:_��1�[%����6�E}��Vv>�y?-c�|W���6�3����z���������6meh*��ķ+��f(�hi	���f�v9�Y^��Bj��+��E�>�g�	�@�.�5�MS�B�xl���� ?45}R� Ӑn#�]�_��+�/��?c^��V��y��9J'��`4]���G����C����f�KC�x��ν�Q�}_[-��F�(�6�;$� Е�q��_rok3T����P�ᛶSc�(�0���z�7����-�ݯ�.�o̮l6qҵ��T��B������8���pK��{��3gy�d��)�N��\�ޟps[�����'�*D�K�B`w��9���]�1/��@�aE:�<w 肷�E�]Czt�KUkR��c��J+6�������I��!4Dp�@�+�a�1S@�2��LHs_�#g������N�>/�E�U��v��C�oF��B�뀡��K'�}뢄9���, <�fK<G���>�$��~�n���ܲS�/�ɽQ��!���H;-�u�a�PI�M��1)�Q��8e�Z�/K,HkU����:�`P�B뮹�u�R�Ȯ�L͗���(2a7���C%��9W��M�#A䙅o�h)�L�p\mi���jڈ���\ ;C�"��T�A���"f�k�7���/,u���?�l�x�Ƞ��B�4
�M�D��>��l�>|'�^�D|��Wњ�"A"��4��P
�&q6~ '�y�;�0xQ�S>]�i0d��˺�f�8G�wK��N�B:w� ň?�y�-��ql{ȉ���̇~\X3�}��l�^��+�c�dթ��f���K-y܎x�����ؕ�����)�K�4d`�����b-��豔�݀獷����ȯe(���F�ʭ�Z#�vk�V�L+��3~d�@�+���|�L��c��]Ǎ��Y�=\k�iV��j:ІBz��ʕ��z��Rڅ�٪L�յr��?�n�YU����:������rF��#��8�f܃�P���A>�h74?odcV��+����������wS��6X7
������,�������w����.F7�f�/��xo�CHIn/��{�����������*^�cۓQ�����i�{vz�,�~�5g��z)gu�;���[e���Y�_�TxG��S7Ef�<� r���i~�F�$��ګ�A�[.?�y鱑�9>�ͅ�r�&En�cpQ�q)�����Rb�jN˦��`��e�i��q}ghF�{��v:0���f��Y�I��
O�u���RE�L���9h����K>�v��V�
�!��:�_j��̮˶�,��K2w��'�Y��THq-�㔸�����*6C��)�Oxւ�b`J2:�W��,w�����݀���T�យ����+�1���=:O���HF|��f�_s7|J�H��b3����DSx�2�y��4v"��(�Tda�'K��<.����ʐ԰����0YM�!R�+��ꙮ�KVh��Q��wƄJ5O��T4�Kؑ�yr/�O�(���t�<Dw�mA6�k��(lN��͗Iy��E�ߓ(E���E=zI5b�0��3Ay����ʕ��2#h��,�A �2����f��RJ���%P���X��w;y����>ӥn��w]Gf�^�}�BK�&�����V��q��A)���#���ex����ZI=�ą,R�����oDɹ�ib�K�E#��x��eJ�I��I�f�c�J[�Ċ��lL"ڙ��<	< F���Q��1ʶ�li'JCWCf��wUeр��`Qc|�iU���N�[){�x1Q���F���K��=�1�>	��p�HE*�rne⢝��S�.IN�ʼ���V�0�7��$D�-d^����7�M�li6"~YV$ j���M� .z��A����~ �����e�j���_O��� ����|'���VYj�-`(<#��Uj�[���z�{����W�w��5�#M��G]�&<�zG��X}[O�Pd��6�@�� 4��UA�0e��Y�W� �.r@��i$�[Ec�v&�x;{4tJ$�k�u)�p���w��}R�f�Y,����Ŵ�Yϥ	�	� ֩ej_��n*��?����LH�7�^x_&>�7��.=g����JwkBk'z�M�ί�@	`�W���u�gjsю��!L�D�M�SWpX�0R��Ŋ����COB|T{�GL9��DЦu;���9��&��G����S�~i�/`��#x�Ȱ��H���
�)�0(�T}��Zz�q@s�=X�sw@
7��"�r��7��n� ``�x$����<$.���]bMʌ�5�3��\{W_�l��%.<��%�Wf"rb'zU�d�O�T" @�:~l�<�p�D��x��
&�]��u�C3�oD�Qo��E�����p��H�|P�vt;���b���ĵ�Qvx�fx\s���@�j��I��@z���i-�����)�\�l�ܰs��ORS)��J�{˛��+A@1e'6��á���f�� cO14X�����2���4��R2��G!��]�_�y�����! ��p�)D�^Y�e�r>&,��5d�l���68����p+9VRR��XkU���Ɲ�+8��+9�P����z��\U��U�)�މ�+���[�+G\l�Cलۊ� �Z��l����a)�C�������R&���x"q�T���,�~�3�%�4���U4l�m�(�������BIFMч(Te�@/ 8�c��>�2L�U����l*�n�!�N��n���)������!��3�f%��W�������pk3U�8l�<dmș�~o�l3��Jֽ��i��"�X��*d �k���D�:�*��2�����,A/Q�!j�d��gI���� f�DГJ�����GIi����ᦰ��bx�CpdqV���F J�#b�4?�=���S�@u9�D.�ڊV+/4�p=pd�sJZCF��Ǆ�袃�tB���v
o��%���G���0�r���t9��L;?�ٟ�����N}���,ϭnƪBƶ���vZ_W�i@�����켌F����IL!` ��؅���IXQ)�Z��ݲ Y��K��Iw�����UG��������ن	�kl�ę�l�\�4��qk%T���Z��zS�Z�Q�C����$�s��<]�o&ޅ�N��܅@;��@a\T��JuF�����_�5�e������k�y��B�U$��!0 vw7<�L��}DY�(	��T`��z(D�0����GD������yۈ�?Kԩ�Gn/��IKKZo��Tߠ���e�a��_x3�q�-[�QV�5(��h�Z��.-���LZ��^E���1x'"L�aN�T�~\�E��:��'�p����
	i���$��j�B�+p�G���~5�[��uЄg�|]]�w�EgM��� �k&�U��肓u(PV���72؊F��k/sI��;L��o�>�ʰb���j�,k��#|���f���R8Y�M���ھ���!&2 ��UI�<�{�5`y�ǈ}���P���T�&��ׇzh�+�~�t�� S`A�/�P��#@��F]�ZD��Ӻ|&}A�`s�������Y�ͭI  "�.�9@ŭ5�vw��]H�_�P`����xL4>Y�lFZ@h�\��g`���RH� �%�Pn��Sj+�^;���	tJ�^ں*�?�R����Ub�,% F�Lj�4a���L��ι�z��W=W@�C2Ű�ƣ�KxD�U;��:Hf_��Z��@�7`�,�>��8�-��{J�ee��I�5���u,�d��W���,���L���J�	(��]���	
)?���Zj�{����Ln�"�־/���W/<�^"<���	ʰg,���>77�ȉ9l�Q����w4�,�Sd��C6^�Z ��
��>}�;B����57P�y��6��3�����ԭ�F�������׾_�@F�{j�'�\���c4#rlA�*�����Ly+��ԝ�6]t�+���~P���y��_�v6��&�+�ҳu d�Y���m�Qbl�hD�'1=����$� �z�t���|08P��PF���`���Os��9�p���zS��]!��&6����'i���Ҷ*�� S�¸�QG��Q���]���dq!v�>�U* �f�X�KN�C�L�-�Pc�Rws�'Am�I�|>,�i
LƼ���}~k�������/�OG��V�e��=����U���w��K�%6{l|AE�s���PRO%Cg��x�m���ر]0]���K����'F�����y�r�bLA�����|��-�d�V�2_0hqįV�MJ�O�`�^W�AR��|\�q�B�8t)	)�E���Kh=�ȦlL�!�aO����h?��݂#PgG�8�@6g�3��[1"�Q��\̹9��Z��� 4f�<P|&71��kx%�1���$�)tz=��̸.Dn
}�}�;c�Jx@(�,������"�u��W�O���+wF���$x x�<{�k��ř.�����S�����K��l�� ~WQ�\�L�ޓv��\ �q%��,sx���AD$f?����؉Qx��R	�3�'�~�'����=��0,/���S���MF��-�������̩���8�("�幩M�7t7���K��e�s�-�q?���Rq�)�Պy���j��<c�Y1�G������ �9������)#U�-Ԅ������|�GG)j\[��o�MI4����������1����A"\��u�[P�7�����NRtE�#Nơ)�`�Y7��$S���������y;��-
���O8�G���;���28?��א���&�����2.��B�EP#���\��� *���g���<HDA������B��r��f��>��ہ،x�$��0F�f����U�ث^)�~~[Y�I��-�����_S�#
�߿��ߗ��E2�5B˽��KpA"@i}��^��C�,�>�g��K�tҫ�&��p�	1gD؀���,�������<��������ۯ�q�
K6nx	�tk�x�ٝ�T|Jiͅ�p�e��8��jAl4��kս�2��P�C��BbK�->���a��T&�$;�i������?��y�S�L͘`%������c
VA"G|:���.��R�����2��#bR����B�� .ؕ/� 	�~�ؗ��5VAvSPB��A��U��ڔ�&
?�'7�+�:�<x�GB��:Cځ񃼋KA:Pgua��9�`��3J[Ys�?�oP�@�9�5��l��Tӹf.f8�f#:�������/ց��ZC��'����z�?QG��({}�0�)d�	1��Y�Oğ4����U^
	vj
LwS�U���b˺r�8�J�����R�q�����a�H��OlC����'ڳ�	���2A��/����d[5�@|ӱ-�q,���������q5�6<���"���zr�-��l�55�nz�=m*�`:,QHpS��,��dNR��[i�Ow.C���6�A�0V�ZP�IX�A��J9��w�R"�܉���� y�3D�x���k�*��mC!���nU#�D))+踤���P)��q�z�QK��[O��H�Ax�� N���Bs��a�g��Q��9�-����#�$j�a��ӀF,�tL��A0�����Ӥ����{/&���EI��3��3�
���3kk�1c��h�	j���i���2WR�m��O�8p��L�Fj��I�`�2"V��T��Q@���_�}ǀ�?��:s6i�^Q�^����|5;0���h͕���Q�l;�� ��ș=QS[Y5�
��_�������2
 R{�K}qIiK������ƴ^�Hb�0 5=�z̄�&2|�W�yWNcY�%��q��Q�����8e���پ�?x�O4>)�T�8�Hf7�U���xS�ިC�'�ó���]��C߭�Y�ߏ��J�c��#`+�6}A��9��J���h'��گ��ep�A~[�p�<���nQ�!&��U}�Go��c�	�a�q�3P4��J����Ô��i�.o�e�I����K v��,�����Q"p�g\a�'�js�T�{1Ln��i0)۫Y�yS侁%��c����H8-[�����OH��z�R��K��I�͡�"e��t�c�l�Tw��k�gU��v��gX����{�k����Z`�A�����c��5�PChP�{"��E���{�Y2m;>����k
E�<�T�d517�B�2�� ��q���p�X�� mP#[`�����%;����ꎊdh�D��'v�/����������mi��M8?� !k�"��Bd�:Rt�(���S�A�@{���:We�������L~p�2Gx�5������.\Z��7:����U������[��h�Å�,� l�q���^f^^�}E��wG��=#򸄭[�	`�u� ��9am_��=�%>E7L6F}r�Q�� s=K��E���cpZ,wH�J��J��bu`ٚ�a�ŏ�����X>�+� �ݸ��],z��G�#F�����)�ς�O9ӿ1�+�բ)p���f��}�C@�hH�kp�w�!@�������a�g4!���e5�®s���Cs?,�������L���z2����k=��:���&P�$ʽ�8�{���N�ˣ ���ĻD1��#Ø q���%q��vx��XL���&+S���-���%�����&ǣ�on�,�u��O����Ά�[��ʃ�-�ҵX��|n�R���Ҥ��Ǭ�.��aϰd{���n�	W����t]�+��ʾ�h#�����G��A׼�)�~&)��Zya����J�;�wi[�5�z�P|�c�B��5��9*]�[����Q]bh���P$�}�>�0D�*.ʖIa��G��(�3{��,����46���n���|�}I�#�k�U�@G��X>&y����Y�/Ƈ�b7�y��2����\p�`��x( i8�)���"(��G�F���L�f+�Tr9�pM�h	h4b#�'4ۘ�+0K�6�ˌb�T���Qv���.(�?2����B3jy�;x��et5�J�:\���NSR�W�߉n�C�6��! �%��&��iX"��I�h�I��U^�����0&,C�� �a�9,1�mAP~������WL?���;3�������~<i�,���{�n�|��j�۶��"�Ɓ���^�� 2��g���<? F��l4��g��4ⓛh�%|j}P�I�DG��������m��t�d�	�X�5�`!m*���uL�?[!�^)���h�mU0�=b��b�55_�G[P���͐Dgz���8��&�c����Xx�XAsr�=���Ņ����6�v�O��E���q2.���S��ژ�ە+�w��*��Z�ᩩ>��lzQ�V�B�6��r���p�P0ԣ�`�6�Wn�bv*h�g��/]U�a\ ��H����}�Ӧ��! yި�\5�[���$E_fREu;�=%��9��[Q�ʡ ��3R�����l°���8��o���s��FlyԆ#��'�Ir~4�Y�s�u��lh�Y���R�Avxj	�qX�2緙�
�N'G���
�����B9�ª���8{xЊ�Q�t�^Ҫ�k�ҷĳQE>} "*�)�?�Ǫ�����|(|��x���}��y,��n,��-^kC��jD���^Cԕy�SD��R��"m�{7�F�]^�g�XP|!�L�F��|�~Vʸ|��%�6V�1j{�\z�`G��w���7�QG�ڠ+��A+��駞�y��Qδ�Q;�&?3���k�����>T���UA��9^�4��(fN���uw�1r�D"`���	�'i���7�-&L��$�-H���������{�$8!\C��k� ���c�>�o1�Ǘņ��Oe)��xp��Nˑ�7ٲJ5D��Ҽ�Ͷ�vt�B- L �v�=��V$WC9(��t�����Оdf��J!2��L��T���y�1��7:P����JߺSO��x�l��޲E0����Q��#�TP��?�ϥE�?i�s�
A*e����1? �rl��a�)�V� ��c��<�h��IǛ�1�N���v�_��_ResVz�Yj*��>����N"�ۉ8Q�5��u�#!)��"�H0��Ndm�)��/�:B�:���p�^�X����OK:��Y I�"}w���6�C���(	�{�E�� ͝s�9�oNݓZ]^�G���cD�p���ik���dH�m�� �ȶ,ֆ1&�+��+ɘ��Q��P��և4´y���6�sMK�����CȈ��o�:Ў���{Q�+u�����g�E{2��ßI��}z)�/��kQOn�=wQ�&,���s<tkڧg�V�TQ&�~��>�̽(_Ow,���ͭ¥[H"���x٪]��4)��ï.�iF�l���d�p�HK��)�x��c6�q}���	������H�R!N�
�d��i�"�T�i4���и�ED�_�M�W:|�c�ʻ�}tsP�"���Ϡ;X���*��}��Ql�w]���"�(�_��N��{fz����Ƞ �&Bo`[�i�qy��w+ZK��ڤ8���<1���>���h�B�"5q�]��Z`���p���iW܂����>zS�j�w{��g��R��JdΜ4�C)�<�d��^�%��_��a���~��0.��K����/6dO����41��+_�/*���=�u�x *3�B���R��W�kv�a�uy9��q�:P��q�|�`�ڄ߫��^�צH'���8����dF9&����4n:#5\4��/(T�nXG;4��s�yH�� ��ܩ�p���K�(p\��I$�@��f�PF��f�;�T�"\��W	����[w&�K��
i,�/��(a躙L�g�z�.��SQ�)�?�>0�kX�O;*="��x���jY��ъ&�dπYK��.�ƳD�T��I~9�ɀ�
m ��+���CD�q�
�IFl��
Zw�ڝ{7�s�as\���*⒃�������N �A���N�,��nDpɁ �RO@�������

�7����u��V��1�#�2�1���j���݌=��g�2��:�Y%�g�6�k���:��t< !t\E���pq"�Z	eo6Y78?�i�^Bk�4���'Q��`9����Źê��uv��,��tR�/��"�'�}��^��3(�dl��I.�wzϩ�2��!#�dU��v��"Iжr{���h�a�{����+h��5��3Q��� ��)6����[JN�Xɯ�1<�å���>�";wF�Imٳ���W�{ǰ����=N�D�c0�v�����F��f��n�L���6�BW�h��L��y�^�$:�x�%�j5P���8A+r�}� ��P!p��wB��P��7/X�Do�AgH����ǆ�#�%�_�4p�F^��_��K��\�����/�&�Mo����ī0�JizBWy�
vq��V��=���(,K��~J#[ߣ�KUJD�`�T������&W�,�$�98��شy�`�Q{c<*]�}�ȡ<7�1
y�y����*��+=���������T�Ax5����V�&{DK��s8�x�+JR{���ew�#M��v�XS�5�������\��3M��XIs)4���iI=��j��ʻ��,�o��T��y_(��I��?�w01�p֑�F��G2�2g����헏%/���O�;�r�G�|S(��$�Y��)w�J��D/q���ט�h2Xn4Fy5�zd��IXB�T}e9���>_Aד]|f)d]���t�5��罖�ke�m�?+�b�c=OI��P(����i�q������N���F�T-n�R����|?(�����iI�u����Y�/�+zgE���h	�,�����W�R�4��mȋQ�8_�gXZ\�Bu��g�_h+�_����+懰Ȩ�$�D�]aN�ҍCY&	��2P���D��/jR���7��TI]n��%��C�x��*��'a�6�U ���V�}	��=�Pv��������RT+���ʭ�8 ���Мj�qE`������"i���z��w���)��˾}�a!DT�D)_g�FF��4�^~�U��UT�8�q��Epv��"7�>)f@B'�%��ăV�G6���t�~0��e_�ȫ�<�����Q�E^d��U2���h\��صw(]�k��L�;�BRo�s�3����*Q+0s�� n즖�6�q�����8��!z��|�d�M�3|W�V�%��0��k��V2���\����<YI�t�\��vg�Q�'���zM�6XE�9/��`� �ɱ�j����c沎%k�Į��Z�~��*֗4��.L[��a�蟌ů�݆�W�:����%���Q�/R�8�\%5an�x\9)�P�.�C��~�,��G�叮u�J�%��3�Ƒ'ڠ���[�h�����]��5e��Q�9?Ht.\��秕
������ 3)@��H��ܵ��K���+H�ԉ*�x:!���xB�����yA���x���ԺA�A�
�a��x��!:��g5�;~�Z��&�0k*wfH">Y�I�4�pہ@U�/�D��0H�2��T>�r��w�譋r[��k28�g�DϷ�NRSu��k�+�����Ձ:Ţ�4M/��~��:�#D��w��2�ijHg��Xx�	�{�8�?̯��a��7G�m�zM����d���
,~���(�a�������c�0����������&I��D���녶uA��� ��tT��С6d0xwJm߷X!��.[�%C2�fܑ��Y͋�������-0f	���Φu|��Y�_��}���[�X����3�Y��5�h�m����W������o�����N����p�D���������������ĵ�Eh�T�}7����+QY�^f0��eR��������4��)���@M���y�W嵔�%0��|�n�
LJUJ��g�7!�`����2��h>�e����a[��Z���a���������+:�1-,��8��3�k*�Z��rB�����oMUPK�`~����<�
��z~T	dE�H�pR��qȨc2.���a�U��x���t,��H�W��E��?H�7^Z��q��6��� ��jDD^�(�Q�c��7דԊN�i��پ�'������";�f66Nd�O��#8����;2�H2���%�>�&�q��OX�JK�AL@_�n�Ũ�ر�cI}��y���ѫ^�����
��l�HG>��M]��n�i���Ç����HE�� ��M2z�c"�| �y���}=�'���y�Ӎ��D�iO$UQy{�Ɂt	n������nP �=�����������)5yS�=d���Z+�1��u����+y�}��d�,J�ďHNM��#$�ul�"��-d�cή��3�|5�0 ����Y��X�������[|�ǫBI[IzT��&/a��<C{j�a4�9O둲I}	Yf�ש����/��Խ���CO	�<f�.� �.�
����< .�l�⚮M�(\�e�H|�h�C `@	�1�W��J�d���A�y�����aVu�����7K����YJ�l#?�h��&v��K�ܯ�����6q���`��F��8�� nl�-w��`H�����ph�,wDf+��k�e�6j��$����N5�K�m���;'[�E1�����:^��_O|��҃��(�$u�t�Gjֈ�v��X�L�/��9�M�h�e6�ÑBX��{���d�5�n�t}�%�]��3�|��Je"&9�D������9�n�&KһL6*^��*�(���	�������J����މ�0�[3��%���IoC5z�>Ó̵P�j�bU_Qe�ڱ���sT�)��H�Z�Y��4�ZȄ�q8��ӎ���Nݰ;Dw�UDW���Sw�RE%�_5��n�����c�$��-����<!�&���Y~�~�h1=���7�Mu�I{ؙ,��n�u�Kd���;���N���}�@:�=��N�nm���������#�>�Fgm�ب���b�*ݞkA@2���r=FE4T�_�Lz��ˤ@��� �Q)�҄q�a�[2�щ�����*�~� �L���V�Nb8�����)�Z��QWvA�4o��`~}�lM��]�Fb� ~�����>S��;�u�?>\!ϕ��E�ET8���DH
�5sU�Xpl��*4[RB��1^�vW@�ySJ�?�ď1Ϗ��+�┠�����p�W�+�!
?o s�?���:�V���>��q��@��BνE�h�ބ��J����5��,��� 2j�o�euUH6���MZ0]a��D=�����S�o�.�m�hr�g�T���	-��y�Z���FP7�������ܻ�B�US�VJ�&5�I���C������iha�M�K-��S�,g���L6"b+�<U���my)�`�頬�SeN�)�7O�M��պ��ʾ�/�Ha�K:��EkYS��}d�$~�fo�N��W��!�4M����8g�i]ӌ�c6�#D��� HV��r+�+5�i�ָI�?�=q�A��&�lj &H�=�OvA��9Z�̚O��� w-y^�����9�E$����P�Dw:�*U
W��]�n-�{�{�G��2p�`JA�5�<Z��Z��6�y��6OmH1�� QRs�g}���L�`�W�E�ɷFzj���M �Ϟ��x��&��c���u�H2�\I���	�$�b%\U;�Lp�U
�b��~֜���3��'���VL~m�4J�ߋ��{n����ݳ$��̬�w�K�{ �P]�4;���[�5��`l�N.�*�����H� Րڇ�!����/p�Z�UK>%% U��]M&�1��j�[3��t�vkcN��y��NI{�ȼ��?��AT[D�]�裒l:�҉}�Rk��������%zlY7��{��`�(F5Ǫ]��zX��9�3~�^ɩ��E{nDDe�`�������N����l����pX�IQ���߰ZJ�u����=A�ɹ��N��j�C��}��U�]���+$�5�fн�#~S)y�SI�kw������by>����,i��;*O�$��L���%���i}��Ȝ����HJ��7������� 4���]aц̤Bc~�;{�i
A^��BQN=�2'O��%���4�5H�E!c�63\�׻�� a���cKpE0k���r_�E�p��3�v��ӓ�}��^P���gN�c�y�J,�g`-V!M��ؚ�:�!9�-e��{��	�͖�Q�׷.u�(���S�N�J�+}١��"Q^@upZ�wO5����w�@Z}�
k�]z����%j���R�g��q���&uf�����������g��%D\�� ��C���J�d�N���6�"�K\|I��R<����!��9�����Ky�"�]��A�hk=�)9���,�Ŝ�����l�݆�ۺ����q����>i�~`��r{�|���q���Y��r��4�f8C4A�Ei�H��G�a���&��}p����A�*�?�edv�n��1)?-B3ixs��@&s�=��3c�k�&�y���r)}��#�x�^�N�ώ?�Sl�Q������SÛ��,n�)�T�vb���,�cͲ@$b)�v'��
��R8V�=�9F�;9s��c1]/?,�PSm+�*d%�$�XUݹ;��������ʸ�w�.fQ>��j[WQ�TMe���a8�2�%΢�A�Y��'&�",,�"I�������ri��ȴl�ٜ�?B��k��7^H<$>���F��g�l�P�6�q����J��0$D�K�,���_府+��%$��qϦs��Y��[?bۜ?�6��kV({.�:x�����w3�v��a �"��-8�O{����,l'E^�YB%e@x���v=�<߰��t^��dݯ��~�ՈZ� �H���UH�77�o�ǠI���w�*y���\}�{�l&u�㚅<-k�~��03Jk�h�/=�>�т��S5l�8�e��\OΔMs@��n�(r�2K��]��}z�~���]�fKX_W߫ b�^��A��:�����3�Q"�|��јc�N�u\,}8Wgoz��|��\�9N�P����L{w$��)d$�p#d���w��v��L��p�$!X�M�Y���.��J7���#��P��Z3Q>���g�;�ꈷ�Z]
��ʀ���Jn���Mj 1�4U�@j�H$�ԏ���G�k�6�,�s��ç�u	˸ù�܍t+� �����i��� �@�/:,M��ֱ�N����9�w����E� ��SQDŐ�I����g�E���¤�Eu	Ov{H�Qr͚��jt ぼ�Z����}IP�΁�g�£K*j���ޫ�&�wO5��ck\���&#@���Cӡp����ξ������i|_�/g��w+L������a:�]!E�Q��l�c�Y4���I�<P6r�#��8��ȸ���0��{ʒ�9=����q����P���h�
���a�N6Mֆ��@z4=l��N!�u|!z:,1k�$X*4�"��Χ�1�z��Q�vG���`b��D��ߥ��B�����YJ�V��K���Cf�/��K�� J��g�b�cun=�Ε"?�P�j�Vg㇟��{�8����>�ȃy��W��L����i�pP����I@�f>qp\m
x�����gf���[�C�@�����%~���6]���b��ҥ���*#��1�c�"cd̾�Ӵ5�:���88���=�*d��W6
~�m�%cyƑ�8t�{�{�<�57ƹ0����cȿ+{ĸJYb��V:�W�J���t��X����A$E|vx����Co6%�L˲�� U�>��6Y\Y��_�"�/�9�4�93����|�)�5�
0U�;T��5a�6AH�4���-�\@��S�	�ȧ.5�b쪭0�kԉ��I&y��i�G��-���BSZK��6��A*��`3�h�dh���X����(�c?�,_@�#�7쾐1�L�ũ�l����h9��&�+"{o�˾�=߳�����jʗ)��{��8�ج�/u���K�� �*%O�Ν/����0R���w�������.��]�˽�}
Ȁ����/�ݙ��P�۩W�j�u�~z����e�^���f&gl�y��a,%NF�H��)l����q�e�jb+��^���ʆE�RoD��'S[-�>�H�+��>ق~��Iύz�j���G�ä�zY,�Y�j�W�4��(�Ԏ�4�~"�@Z֬�,SX��yc�k�w*c	��VGI|���<]��#�/��-�#]?���{
 `��s[��Y,��ѻ�qjDW�}��<���b�B҃��Z�	����e��E+M)p��H�b�hm�+t$��V�d�q��:��M�Z��4�ln"W�j����/���ZJ\�6C�yRe�['��Lj_@���*��T�(=��aoA[]S;@���2�d­�V]��t�D��v���m|�����L�0?41�h{-ƺj��^}�;����^9�<��8^��b�0����:0Ip��E�2�	�_�rwM9���/u/�k�5��oM�?v�UԼ��no�-7����fU�����ᖐD͚�:���:锾�	Iɭ����ҷBz��9d��f����_4:�ↆ�1���[΢��\*�i���e)QO=��!����3�w:ɔ���>��aU0 C5{�m��+�A�g`Z���q`9����Ӑy�R�Һ2&):k"�����d�ܿ���D�(�c���x���O�u���w�Hj����sמ'Q�3����8*ßű���Fn{HN��������F�"�;�=��Tkc��wk	���$3>�������^��X��Q��`�B���������*(�4/l) ��4��@�w� ��c\u`�������wfU|m��4$?��yX=.��ǷsZUF��.�r�R�=���2 ~��Fܚ|�,�CBGd��Yg��eV�9��s�q�<�N�E UԽ*����;GՈ��
']~��!��Ua�W���+:�Dv��(� �,������~�a�H�̢�q�����w*�!X��+9��/��lX`�ヴ�oRޟ�k�D�d���U�KB��+��"B9j�N�f�⩑n ?6U�4��6�R������&lsp.�\0��Ep�RB:�vl�M�ȕ{9�c��Y#b�+��� $�}�d�M�q��'�ru�zF���
:.uyX}X��a~+�kto�!�
��i�����}ñ#&�Ųթ|^B#�@�\��em��&иO"�S���(�ъw������rS۝����m���^\��R�'B���h3BW�%(�D����ԧ�Ǻ"p�׽�'q���h��4�x���F:�����w�cߞ�,r��s�����7ҽ�Xx8�8�t�T��� ��Q��3�++�LB�X(,�{7I^��9����} �J��<��q���q�zǜ�N/�Ô��(�L0 �Ԋx`��@�ݛ궱"r�EAߍ��/���t�ߐk˲CL�y, K��&�l��#�u#�.�r��Ԉ1D��OO�����[4Lj�A'�\dߝr�O�ࠔ���/���W�ޤ��u~9D_o��A�,�Ru�ߊ2�7���f�1��$��b�&k/�F4��tx�����26Z��A����2I�����/��g�(a~�^kb�4��ܐ����`�s�않9�1sn��)D��X��ǖQ�P�$���J
:���_�)��pW?� х}]:(U͎�{/.ཋ/#-`Gj��Uzo�CF��n�~��k�~ee,������)@9�g"䑿����)o�x�|�I�����t:]b:�k�	�z�G�*8��ys�/l�Ħ�c)�a����a*��;$QuQ����0cr;i�q'�,�<��y�A�!������ȸ�vCU3aZam�Љ�/�ޑ��(��G��)�3��eU$� �"�:�-�3*�t!����1��|��6�'R��U��3ڣp��=���d�,�G����ޥZ���-�͞�^0:
,c�������h$CR����f'"�X
$#T XvTú��|�6����b�\�ΕVW��5ܕw/�ǯ"���W�_I����  ��y����<M=�����M�C+��	��8�.U���y�ZnK<e�G��VַW*��.����_ijz,�P~�ʌ���.r���Q><�J���f��0.�鈝�6`x���!Uy ��0/ڢi����2�{p(�o}�Y$�Ȑ�rםnU�l��x�[��>����K�"�j/��q�1���Q�J�q1�9Q���g���w�� N��~��B[c�"墜P�b��=@r,����!M�8�sɑ��A���9���Ԯ~��󔭛�*w�F�&|�ߦ�v����G!�25x8�|����G�9a��yX�I��7�CA��Ma��.Q��Rso�C�a���$vq	G����XC��l'.�p��%[ĳz���҆V�K����F�;���?n���5g�C" ���K���>®Xry�*/��.ģ���-�{����f
����d�<�'E��B�M��"ya�H=�@��qg6�3�Y���������X�Xʋ"��$��}�{��w�(��E���#�GH����d��9ȳ1�G�����"Σ~2��R�뽰F:B�L"�7�RbX�QV9��Y�ּ��d�Z�d�.��T��%w�g#�!�0fp���e��"� Ջ��7泗�R�R�|t�q+y����*�n�M��d�V"7�Rm���X@[۩�fJ�8Sg�15�'���0(�xE����P��}�����H��2����v'�G�Q&Y�yjr/M��y������s�������:-bPT�[|`�|���o��H?�]H�m�qJ*(�`�(��2Q��؄��b�n�Ka&��'H2p_�	2�y�|�����F��;ȋ��v�[�g.���&��+�Sp]�	�w~Y)�v�p��w��*A�;ݣ,�Fc����5�'xl`�;�J5@%�v�����?8�+�&�O\�SMN��%x�0�dmܨo��8���^F�O��t5��.����_�m �x�e��E߽N_��4�����/oGM��ۼ�`E���H��ʏ1O^j�^{Z=�Pb�H=Tы�=���y�_=�0���E$3���O�io�F�맴A��9�'�>j�A��=V�}�b%ci��ܛ�|�%$D�-]wIʼmf�x���u����qfa#��t�21�����ί�O��C�`k(�5��<��Ff�y��Ԙ����#b��S�{FxqC�/*�H;��x�#o	�^�nwk�sd!l&��T�֐���"=ю%�`!^k~�ɴ�O!���c\�	3Fm�9�=YӃ��Dk�1��VB6a	���FH��QU4\B��f͐S�;v�N"�}e��ӊ�OEU
�J".���Dys��\��A��ݥ�m� Ⱦ��$.�t@�:OE2���֢��P��H�uޒ+�,�Vn���C
��s�z� }�87~$���jȫf���р:=�@���@g����>��G&�C��H���
۽{-o�P��I;[O��D��.�ҡ�y��U找BO+ZL�r�n�`�X7��XSFm�{���Q��Z\��`�u�Nd�k�cW`H�K�)CO���Ny�*I]���<B�.���mC�zfV#z���d��B��e���� �q��Ùagm?�!���2�����IS <���ar
����߰f6VF��Ĉ��sT,�B����/^]t��%(+M����}c	�.���Z���^�R���mt=���$��+q�������[��,�O���-c�2�N$k���6)�����Ch
���}j���Vl�����������U�cK�A�L����[�։b6�~$j�u��Ej��ίh�$X����"�0�Tl�6Y��V��^��\I˜#C�}�6 �H9��v�рc����^��~�*M���X�*��[}�2�9q�RN-�J� �Fn� �ƉV���G��4�;�}��a4�F�fp߂�p�Ɠ9�����J���V�oK
�P�ɸ�m?����X�6-�-�ޯm1���>�r��a���.��%}	��!& I��t[����,�U9BH1H�v��X+��P ����7��:��U宊�|�<j�{sc�&�e8م^����%�	�S+�bdW���F����t��7Uߛ��Ʉ��7xo�fp�$[û��.׹�H죀���v�W�����MDƮ������q���~�Mm
�jJ�e&P���m�x����L�tS[Q���W;�G��	�Y�'�@Y�����/��)G��=Q/��C��
��!���+�C�/^��- k����XU"�Ɔ���>��kt�V��`O@N�����+��:w�:��I�q�J�Q�<3�����V�şD���BL4b{,�u6C�:�����N$@���]�/�x�ǆ:��Bd�5��-J@��Zf���v~L��!@|)Ǭ��� ʻ���*?�O��q�L>�B&���>r����Y���d�_�'Ǒ�'�T�7�v_洤����}�ܓ\��e�?#��k<H��kdZ��,��UL(�6#>�H伏v�:�D���22�Ub�f�TG��g�����*��Q���U�M!Dq�'�i�*����]Xڵ_��O�-�����G&%�]-��2��|K5�9]��������Г��d��m@_�K����-��8��v]LqRV'�7���5p/��w���M7���2��P����؈	�,c
sD��5��<� �� ;W�P4��sI��I���$e��ڃ��œhd�?7n���a����x`TJ�,��n�yͶ�����nJ�R�2o(�4M��eⴖ;��\z°�~��a=�ґ���j� !x��"�С,: ���{Z΄G�߶��{�΀=��I�S�z@�o�����ҳh�`}�R�/�o��(Ï՛����������Fa{*��B�=w�h�.��aR�fiU&��V�5�n���m��E�]����`�t��y~���x�#�W��/{+��Q������� N�����̢r-��պ#����3,;�!蔢�K6۳W�]W�QZ��1� ���H����R �TXF��Zʽ�x
���z;�Jfz���7l}?p����q�Q{�f�vfPU�	6	f�[cE:��>���_tW���kB�.��]w�1�Y�_E>�Qd��z��b�i_|��a�2�.�e�̕��$�8o� ���stMz]/j���{w�]�\�`c�x�RO�[H�� }���]fU�]�du6�����BJ�1��`�}Vo7b�� �p��1-�J�d�EjBZ_�q�F~.�4�p����x2t=�Î�1:$F��K����'y��Jt�A��ߵe�",I���L\iLeL�/6�M5�qe:�e}�5��&g��>����0%�����Pы+�oG� 	^t�D8�ã K��s�:�L�q+�sQ�ڡ���v��%�*�㡗0����u��-�f>�0a�2�VA�q۠���IM����Qg�������}��k2P8��������/`��w����:��EV��n��o;�����򈔁�7-��$C���%C�:9���Z	�0��9�o��G�
�[����yt��^��aK�A����(��P[��&��=�պ�J���0�f��u��hy��h�.4sG��X�t}���Qf�@@��R�ERU	G����Wc��9�����s	;wy�)֬5��O*�F��0�1��2~��<��Y�@��M�6�)T}y�,���c�P�w���O`!�>�N浥���}Iq	P*"�"���U�b<)�w�pf��N�{c��rL�tf�#-6�w2gpIL��=*x���:R ��8�O��L��(�2(rc��P����8�~�?�|�,���@iV�f:�rq����c/��~������I�u]� n7��|I��ܸWX|�U�>���<F�|�v���2��{�� �Y���W�đm��
4��{�yO�E������|"����,TD[S�Ǽ��jv�5�i�S�BÅ���M̽�����D����(�E.��(ߔD1�Y�t�׸x8�i�h��Wn�@'�ԥ�gl�+o�wgDR�:z>�lݎ�h�?e5RЪK��q+�5��Yr���a�ؼ��M��{ۈ�I�GOs�MW�~kǒ|d�4��S؂v��ײ���� �/��f��ji�g�u�ѕ��3��x��G)���P^
)�r]�2Ҝ5���B)�U @Q���֐��I���w[�*�'��Uqj�V\�0>F#K��Q\�i�l�Yg��Aɾ5���h��%�|�S)S�Kl�>�� ������F}��Σn���<���z�R�G�4��}�|�.�3'��V�q9�M|e�Nj[�� ��t\t�T/C�s#��d��d�y|�2�٬X�ˁ��#m3��V���{��'�{������4;1T*����~(98Ab��349�t�-Pn�|*��bO��`RrBO�K0���*����:�K�uK`)�y�/��|�n��xL��l���3o�f�� ��w`M+m���0����r cH�͹ʒ*m�zΑ���jyM�Ӡ7R����N�q��h���'/3��ԑ݄��� �cUrdt�JQ�E"W����d'.Dd�v*h*�JRO|��T��B�E��+��X�2��F�9FۨXX�o��%��n����C8yR�s����x��C ��EUhx���"b��Ţ�_�ܐ�j�0Թ��t�Z�ϮG��O�k�
����A����O�PGR'BS�v��'&A�Ҩ��kj��Q^X"�:)�O�����D*�#D4��7%�T:���Y]��x݄.�Ԏq�����7p��\̓n�%OD �7�7�w�ԃ��3���Ёx����F �}\�l�*f:Z�������n�M�D�(��u'ǣY��y<�/�Y�0y-A7�'5��V{}�ϊ;_O�c25��������@�K|!��
^ub1�d�Ň9����b���8D%�lp���wx&Le��v7^#���;���I��m�#�y�\,y���HW_\)l2MwKt#���Vx����-�*��˦[6T��Ti�}�Ⱦ-5.o��S�mi�y(*�xmz6�k4]�hOݢOL���J�p��d~�Dv���/�R%��\���&N�V�8�X��ޗ��;�U���|14���c��C����ོa��^|��>Y�p8�@�ЫX�]�|�.B�B蜅פ"q�t0���E�0I�v)'/
^~�?V֯��'=W!�X܈4���%>����n*](��E��X��<﹫]p��pO��_j��7u�ѭ� �*-ԡy�mq�z4B�h^+��d�#�>d�F���i1�!ś������(��<��@7j��Jx7r��
�8V�4svӆ�$iV��1I�K�EUִk��MYx��>϶-����?U}5tPΘ:l�Ł@��<���՝�!�_$#��j��٢�U	k�7�|Z m�����cm�6��I�nq*	��w�h�gd�^�(';O�.������:6�r�OP6:ǁ�^��]Tp�*	�u7�r��a�M��1�V7�X艆�E3YN+V�������?O��e���\d­�ߊ+�2�_�?	��#�s6D3��%���-��zߣ��j�n�E���c���R-d��u��`L6�����<4ہ�];�Pl&��{E�\Od��_U��]����Ϙ֫���Q�����XoGsrU�4�U�c�K�Ր�M�����ϕ��g���2�4�ڼ��R)S ��u���Z���2�NF��f�	��t����=�m��Q�)���y����Q���K�"�-��ZINE-Y�K���q�+W��s��E�'��	�sv'p6�!#�R*s�*�n�ٶ�[���U�s��O&�X��<ИMV����������mv�$��r\�>H�]䓓�
�5���v;	U��%�� ���-M�	G�7��,@�r��)C�lA��䨯�3��l\\�a2�l�b���0����ir���}��W�p��1��3L�`�L�?�f6x�dv(�鐥��Q(T�q �|�)ٸ�Q�Tp�+�g V�Uu���_Ձ��ǣ�3H��,���Bu`��4sͶ8V�d]wC3��+�6��X� ���{����(��K�xf�ILW� �}��2b��n�����	�Z��b�o�,���LT��T�0@��I֧' ���h$��z�s3YQ�N�O��D��(և�=�)����8.��I܈K�Z|��X=E��<5�c�2������S�ǵ�ɛ�� �GS>�� ���õ��8�bh���!��:]p�_��T&��
}�K6�Ym�x�_a�Y>�@M�+�C�a�{��7M�v�����6~���Y�� �n�@촡��JК�8����B��v�սR�����?K�����p�AD��x�D��{	���i�M+j�g�:"�M��Ӓ�±+������G|vX��-z�F�a�ҷ��1ۍ�e��=���eOڌ�.Q���7s�������1J�|�PG�q��9�zZ�����!���X��vɒ� �z[8c�ǽ�lKOq%c�Bfj-�t2@G5ٰ�с��E�8+���6��28�@�:����v+��:���8�P͙ ���&�7w�O��.���x:���^���7����l����Q�J�򦦥�u�wc֮�>�	��'�t�Ɵ���c�OCL� �82 s/]�p&F�:�	���i��~5��t�^� #��iw�I���9K�>\	C��gw���6]�?s|�qm�܃}8�M�<��SƤ���7E=�$���w���vq0^�]Z�x?̾�d�I�[1�HY�\�H� ��8?bTN�K�j˹\��-����&��8�S�,$���t�y��r�ȋ�A����ı-���z5(�R��5�\�ָ	�E�pl�I�gfrBM�߉̠��TW�2Ӯ�zq�uH��)�$ �^%�ރR�d:��ِ;�������Ù��� �d{R�}d�ة��Ő&m��^� �	��m~)}�6����"c�L��i+jپX�|��_�X��֣����� r�;�r1�xp���M?*}�%��t���_fwq	���+L�0��yy�_��h�/��I�]�ۃ/,0+'�U��H�ZV
���N���} y���r�훙�'�	���n����V��׀ ��9�(͉�P�����§��{@���C$[`��q4�6���AQ����kS���.���2�����'WQ�`�z��_��*8��0JnX�@"�\��su3 �@]��{�=���5g�Qz�O�m<R��C��n}����߻�N8�����7��p�&d$R�PČ��b
$� ����T�;��(4 4r��۠ș�HP̾p�I��_�������33<����Zy��<>���K�Y�'��W3$!���N�z�S��:��b�l:��3��㨽����N��ީ��V�k�S!:;��MӒ�;U�e�8V�Lܬr�	�)�h�|����J�N��_�g��8g��/���C�w�=1gt�Fm�[���	���̞cby����+�B��-�7є��*Лd���vkrhO��O��� %DG4��ZɄ�Bg���
2j�)n�"�H�g?�ָ������<�r��̜�Đ��L��5<r�+�&�6g��6���ֱ?��8JH�[�
�5�E��W��	�6��������\��׻⥪2��n��b��(>j*��0⤿�~�4���.�mYeN�h�!R��co� �O\���C���+r�oj��(_�PO(��d�K��Qz |K�#�o2�K�pJT}N�x~&��'��z��Z��F�C�Om�+-y?�w�I�HN�������(">��2��R��
�ą�� ���n��~�!��Y��f&���$�:ډ"!5�P���5�AW��]-u�v�v��N����i~~<jif��ō��+�~�o��H�I�:@�͞`���;7Ol``[t{�T�+#�-X�d�5E$"���z3]�
�>P�KX����:��٭���na�aX�,����{�׿X�;�b��/�x�M磖>,�ߺA�|�~�ْ�b�m)�u�eo���	Ul ��4� �~�Vq��~���?�P�Sd��Ǹm#�N���`���;�D�(�#k�L]bUɥ�א-�q�Hɓ��^�l��9��+�tL:g����9�����!�%p�7����z&r!_ ��?��׀:����8�r��(��ŤU+��`���6l���2�� :)4
���Q�yZH+����\�h��#�	�Jչ�ވQl\4b���L�1���%5���QxZ[}�e��9^���!6x-<���c��t�4İ�\�W�̨�l}nPz�8����<�ۄ����<R-j��;���r��^tA�3IFM�.#��:��W����JD�k����F�ʍ���	�Z�s�z�x<ظ��%��;l�u�	&S�1�2^���7�~?M+0� ��:+��lĵ��NH���1�!���3�e�����)�(S%���_��x�  ЕU수S�/f;3Q�/��o<{?�4"Cz�'����U@�B�>vz�̼Ӻ�S�B���V܊���l:Ҷ��j՜�����E�? ��	l�u��
�ޡf�$�=S����=���]�$�ԙ��C���_{K1��ψ�ge�-SI��F`����55���tq������6����Nw	��J=_�nˉ/k6N��ʧ�N�Rؼ��+V��Qի�ۭp�)�[�4��!,d13x�}f7�b��Ʀ�!1BH8�qX���/���H�%[����^�ٸ}���$�4a���#�@����5̺İ[%���qW�[��`2L"��=,&�s��+��|��,���!�62b�l��u�
 @���rr��djf51BL�R>�D�����M�8�_�N����9�c�*Ğ�����1A)\��5�/�e,Sx�|�'���s&̭�j�Rn.ˣ�gD���՚+�@9�z�������S�o��(��Q0+�s= �J��N���DVhO�5��C�I��v���	Ν%����=�U�`���F|�s���U�+?g�� ֪�i=g���F�ap��݋/A��^Z<
B�i���	�L���x�5��0����Y�����$r��'TPp9�$��A��k��Q��|!9�l3��Y�< ������H�<n�LK��E���"��<JM���6�qt����=� ����������v�f��FFJ�>��,9��D����>٥��x��-��1��-r)u44;��5>������qBCڶ�=�ytkXq�N��ZJU��f�pE߲®��y�,��s�vl��c��w]�� ]��e[�.�z�ܴ�t{�c���7��������"������9�]��%���WXI��Z9�I�=����꫌k�d��R����~RqLo��/�-�0��.�K43��q>�j�㒖���v����_���Qz%�g
�Q0b1�|�EM>�<�rnO�;o����=���*d!��`���^����V���Ɗ�<�љ-�UkX�m�+�qX������9��l7�v1:`}z4��c#Cb��?.U�6��B�@�b��YJ�Ɉ�N��9!Q<���@i��0h3¯?�	�"?��Ks�nc"����F�#�Â�aW������pDh�jA?5{�25����gӋ=��S�t)g��D�i�V���㆘U�Kgͳ�AF:�$9s�r<G�)�j�c8I�OT2]��}m��"���L+��A�+�%�\`ȧV' �j+��6��hMO�:JT��S���UQ�Rx�*��-@�D�ng�����,>-�4ID��E`W�k ZvCh�89��H�/ڂ�E�+��ֽ�<g]��Qh�D�@�v8�Lh���WY�4��ra_��$��<��h�-��n�-:*9��uB]hVG1AW�q
#�X�dV&�f���@U7J�sSC�����z�'�EPz\��M�n$dtC���7酴����~��������wv?6ݙ�}��Hb�����z��hQ�6�R<U��}�㴹��OZ�@;���n	{�_H�8HR��QZ�2;ݹzp�o
2��_�P��Ko�<Uj1�De:�O:�M/�/	N��A�$�_,|>u��q�NJ���^ ��00��U�)��L�_:�^�_v����"@\UCA�A1�4I�%�G�}�Q6�61I)���h(�Õ΁I��@��Z	)u�A��y�J��XחG���rG��J{�����(�r�XR��t�Hȶ��7ף*i� �$��=(Ɇ���ݘ���N���]y4���ϝ��P����0����M}עU�GG�~6,B�-~���6�?�����lE��\�\�,N���ҕ2���>Ç�;�iXN�U�|1��]��:L��b��d-{�ǿ�c�T?}:�Y,�a��B���Mb�Gm��;{{�"��WeƵ�c��7rqrf+_�k�>F9t�pu&8��ı�$lyh?1ͫ�w���4���z��o��y1y��#aM�E�����-�Ɉ���v+X>|����P]&:���NȗwQNF��� �ݲ�v��&���%�b'FW3?��9���C�k��e��̚b��PB� �U�7*ԙf�8�%\�2�F��6��%��ݭù&
M���a̍���XY�������+��$�%dJ�_��HP�e߿���տ���f&����2%�M*R ���L��;�u{�t.���ϱ�^��{�z@Ŗ������f4�F��D� \�*?����k�@2���s:�鬭f"���������{v��W��^���v�LK���<�qR"�͏��~ZH�[�LK:gR��@��8x��H�=�' ��Ҡ>3�g��A�{h�%~i�(�g������R2G�Bi�H��$��M����Y�0Λ����xmX�j�H@g���1 Fo�ģAě����i�0A.��E�I� �5�2����*��k��N� �)�M(W
t�����F����{N��㚫c����d���N��h��;��	�:O lG�ϽL'��;��<�e��k)�OGl���N�D��d�"��� �Mg,�2���Z��h�cg�Pvx1S�;i9����6Q���]�Tv¥,�*r��z�뼢���5��0Ѥþ+���/��LB[F$y�]��k�����ɤ���ٳ��*�#x��'�:��>_s4�$�����Q�|WO*թ�L+Z�||��YM���($�W��e��B����:Z"k��#@�z�c�^�Ï�+�q�����T��bd�O�&J
`j=���3:ʰ����<�̳��۴1��8r�*����D�k�^}��+����5@v��9�6�-x�򸈐�N�(<��*�Z���bC"np��=}O�㵔���f�R���R7���eк#j�*7���!Uj�g����uC�����'���흲$b��s�)���!���O�����=h���N����!N0���o�e�����q�bRs���vov%���fRs���1�V�s�)����}���!:<�@��I�`� ��9�W:�S��	<��3C˫J|m�*�e��� �GY�ℚ������6&��f�Pwg	���T��1C���c���y��[�*T,~ wNir�G)��0ڮ�.�V��\ΦށԹ�X�5�8>Y�d�J�{���ӫ*��Ғ�X����&��)��ol,c�g#�c]D�}7��X�p��)���I�0Iͪ����,�uB�d��;$>�u�%��i�@p{a=Ӝj>�K�@��ޔ����:����4�%�TXp�S����W7���C�W�~W�f�xR�8��yא���<ꗳ���/!��85�w��m�'�X�0�SU^l�����x ���KR�Ю�Ƿ�j�/��ʨ����E����+ySήA��H���a�}$CT��8+�������M��&7���_ڋ�1�8��ȠAE��p�~z���j)��jE{_-'�:k��uŪ�jA��==��h�%�^�<���� ������oy�M�dUϟ��M�v�x,1}j��yvc��Q���Ca��d
�9Pć���a�|&�k@Z&�0��R���>��'u�����c� �%�>�U?z��]�6�u�������sO��X����FJ5�giF�@Fw���j�/���S�+s���T���v�w
��:���ɒ�!����d޾?Z�SQj05CT�-�$�����bf�̏��7�B:���egah�Ff�ћb#�M<?��p����,�����9��iU�sW�ΐR����	N�xҚ�9UÒ
��r�UF>,=gM���:S�ޠGutS<�^�d9b+
���}C %<�N�}�����t�|K�9�zf�}���b�4��d�e{�#��T.|#z��߂�0�iπ��-�o�#b>�"����KlI#ֈ��D���/�l����.�)U: �N�C����@���D��AC�V3�#�Vr�/�]���ȃ�]�wä%|M\�{�q�� ڶGP����ק�	K�#�f�-轝�uX��h�pd�K�J��Ժ�����h�>�GM�0��x�\�j;��t ��y���2 ��UD�U�.=�Bye���
�[E�"�#�e�a�9,f؇'Џ��Wt��O�R�l���<����8X����v�bH�Vb��*�{��O�QR��>oCB;������V���}���_V~�i����]6� �m�Z>N���� ��S�Y,����)ă��3�,�. ӿ�c-�#�ifߢ����Bw����C���W�J��b���E�Y�<�����]�$��?�f5Ǩ�"�0��D��gʪ�!s5���k��� ��?(91�k̠|���`�P:���ݭ�ʎF��
f%���Y��^X�i���+�TpG�๣�I{�N�'o���K�*Ґ0ȏL����m�I�x�j:��kEY�P�ܻ��Nx�������1@�C��+��ѷ�� ���R�?P�c/�/]�����B~���*���^��8�bm!������7��Ȉ�(�^�Y����Ds��L0#H��* ���3
{d��Ʌ�
�d@�]�4+�B���,�q�Cb]d�����X)�t���g�X>����ZҐ���Fj@��xB��;�A�*�y������V�ʓ�}ՓN@��	yQL>0�(��R־@ ���F���
�jQa[�y` >���Nq����<��}i2�N��j�̰y��y-'�C���%Uef�%.ڌ�C�ȥ�;1��� �y��N��dyy���O��r��j��!h��6���# 1&��L�E��W�2��_V��~Vi@K���q�¥ ��r��ԓSO��o�q���9<9:���s$p�K#&�b ���h�!f��e��ؼY��>���Vr�� � ω�/;od}�ǅ$�d}ˣ#��dCI~���U��[r�,�eKK&yэթ�;�N��d���n�&�u	3}�7�u�EyQ���B~�<�L�� É����Ώ�eb�N�^K;��'�_6��-:k�3��$��e<_T!^Hȕ��^<lV����J��$��L����%]d�6 e�o���
4'�{ܙ��J32�>)M����RA���۰ک5f��VgOvp,��(�y�ϲ[֓����u�,�B�]�K�,o�O�����T��!
0�p�W{���W�8�^~�a�V�z��.�"E�y��P�?W6y6IyO�4�b��<�5�u�ʗ�o~�x<ږ^��h�[l�j^W֪4(b�'E>�4t^U��8��#�.��7�a�7�>�df��L�B����i�qy/����#�Pzp?H�ٶ��약*��'���G����ȇ]>Ğ}O؏�B(�yM_���LZ'���7\�p]��`�y=��C9����p��w��o`3���q�J���PlÜ��G�,�7���2Ľ& ��
}��m1�\,?���W��n[9���r�Ö�񳍜e��|�Mm���Qo�K��W�(�ֶ��,�s���)suP]j�˴��lD.��T��2o&%��݊��Ր���Ĺ� � ~�Z�>�1{��&�%?�ό��{f������n�4��w����t��`�=�0[�r��~6�k�oT��K��E!Ew�s��T�U�hp6+a�C���!��r+��Ж��h���_�=6-X��S��
b�i�8��A�������ő)��Nm9P��'���4�u��x)	5 �E���ľ8������^�'Ɓ�@�TE}aFEX������ -,��Q��:J�w���3��ϝ��ſ�.P�X�����J�
�x�]9G�[��<�5���x�+�uC�DG�j��}�*�鿍g�F!������n��`�\�$���*�:`�\��V�\��F������������dǗT8$��[����ՙ<�w�������]ͤ�W���ZK�y�>�(l��d=�d��:�
-8�@BD�e��>K�d��_��k�%��+>)�
}��(�W_򨄩�m!-��.���c��>nU���Y��>@+���"MZ�;���c�g��yl��"f�(��o�r&M	�6%op���7�ݮj쇕~����ќS'̟��V�]U��E���G�	�ܾ�Ŧ 2�S�/p��t��+�e�{�W�ľ$,}ș]ĵ�Ul%�fX�,8=�0�Q��P}7��E9�	�
O-%��y�R�q��&����lK=d%�M����/��~b�D��ĸ4ADG>����Q�R@�����o�B�H$��q�PW!�7c��m���̓�H��!dED��F���86�Ov8`�ePK�X
2�(|?��z �ԉ}���f��!�G]�*"dn�~ǘM0�3dK��r��uEӉv��7%��1I�xi����,�çƏ�]ʱ���X�f�J��8:P$CU���ȟ�p�>��u��Xꮤ��1��z��<D��i�����;�і�;�{�����R�yiI���5e;J:�C�a���ΫVe�E^����q�1�OߗG���N�K�x㲍��~ Zݍ�N�+T���ohj���Ƒ���� � ��N$\�r v�v	�ث�-�&v�~�����|n��������"����%�PX�9�M�cC��(9�5����$�~v8���T�R���J�-� ���[FD�#����B5�W��b���c1��$=)?nG4�I5�,~,��&��d��E+���7W�P������9��L�[w�ݧ)r;���@X�o�K�gU��+ፖJy;	���I�g��33�8�;j�vg7��@��e�1ê0���Ƽ�Sa�^K|�e� uտ�V�t��/ܗz�َ�%�+fyY���gk�i��dv�/��z�o͂�m������g�{��AO\8���~�`�7QTSazI�D���[̡j��C�ydD
9�"eR�FRt�r�:�_�>���ӧ��F�����nhuݻ��tq���TCjX���y��3���Gp��g(X��x3�a�O޷�����j����O;�އ�|�+'�UH���)_�z#,�>��9�U�I����l�=ٕ�˔���@�UJLWI�2���	����M	���V:�xh%�=�PEN#�.����#�Y�,�<V�*���~����+����qf��
���0t�]�JYhJ�\.�syx#u뜏{N���H�?;�3T�C�Y�5]@p��$��8�2��M��E�s}��Yo����UnT��"�8��b+oLJPTg���H�{႘��h�"&��=/9�Q%��g��,RB������<���)�\�&È��8��؂�Xs�;>�fקq�lR�;�5o�wtCeo_�9�r��xB�K�R��@�"Tt������p4���b���/��3�.C_�$T%��ʺ�k����<V7"�&�/�u���>���#���U���9m1HB�R>���#�g�ȅ"�Ȍ[���D�<��:�O{��e_�ne�.��?e�\XU'�P��vk�yL�B&��0LX�]�q�0y�:�D�2���
Pb/¯U��X�|�T�e�_��\7|�U�O��F�a<ϲ���>��fYv�\�dF^�Ƥ�D�_H,0QaN.��=�[&��%�S�1讬�0=�� ��\�i����J1���#oQ�a�N�-�(�,�ܤ�����KaA0�H拗�����ҏ��=�aQ�*�Sȡ6�Yv�i@�;<����%U�ܴ�o%�H�Q!�>3�*�u�s��*���?�|mҤ<�T���
�:���lq�.R��+yk߉�>�r��R�5��˟�i� �7%�mkY���� 2�2��?-��aV�Pi��|Š��)��7��8B�^��:��W����C8�>쟑C�V��ođ AY����Qs�L�/'�GZص!ؔ�[-dQW�]�}���ۯ����K�`� �Ԙ)�d�NJ>�R�	�aP���T}xA~�p��<w��ѝv$�/�C�ի3�w�H)�G�n.+�d r�p�g"�$U�?r��1ը-���-���cvަ�&wPsz*�J���Mn��?��1�j��t�k��a�вz�׷7�7a�I���6w��.��M�7v{�{'��޼.|�9��0�k+�|�UA'S�"�(��� �w.r�[����Co|[~>H�e>���]m���5_���z��A��BI�x������Wy�dS�����J�'l�o.�{�1�T���JX�������O^�׃����#���-z~��ķ�>znW��i�&�}{��of��#����n(WCK��L�v��:T\�u5�Mw}X ��lM��e��B���n��Z�a�������Ѷ]i����آ1>�\�4� ��)��h�
����.f(��W�KtS�WLbq9�f�3i�89���z�؈��d�6��z8�ם��A�h�'{���b��oLE4:�ԥ��rޫ^z�,��Ϋ �ŏ�&0�������><r�d='r'�q���a�����QEJ�؜��`�5H_?r;��$���k�P��_u�t�	|�"���j��i���t)u���[���Z)�)� ��9���[��u�v���Ev�tp�AF�>U���aT{� ߜ��İ8��x��.�hmʫ:���<n���o�'�h�T�Z��qI�:Q���={�5 �E\Ἦ&4���Au�*fi���$딚����"��=����in�S�{�T���o�)E�\�� Ύ}�q$��iU;E��퐱�g|�
��<nO%��\�_��"�,s��E�ޓ,�Lj%#�`+�9��eD?�7��1c/�������=��Q>�Z�A�f�ao �2@��nVL�� �8by�Cv�1�����׉�g�kf�
�D[��j��Cd^�+p�7����|Ƃv {������T�C�6�O(��S��[Y��`�*���b+&D���-�S%%�� ��؀�?��U�Җ*#�p��1�DGR�(I��� �.��$q9��y�lY�c1kF�W�t07_�Ѡz�'b]��q�Y%j�O6�*0�l���J8�_u��v����y�JJS�rN��:&]�1+S�G.�TJP�k��K�����mQCzvov�]�`��&����6p2H�`����^@�¸iգfN�S�-�^�c��!���<�H�9�5�U�T'{���I�Q���N��;GJ�ҫ4XPd�"��)�W��l�� �8��?^,�����^U�n��B�z%;�����)�D���K�'sM�CF�1z*�K�_�d�Q�>ci�t�4Qd��E�Y�w�f�G���w�in��WUG�>�~��m����������хj�u���=��U�ra^�f�I�Eb���Kl�MzkG��C��/���./_!f-W�E��#�-��AK���*{��Ƙ���W�2���+�١�ܣ!���(6	��v6���E.=�.�2�����)7-�j!<L���Έf�F�g�"����5
��j���ZX�}���s����5��c�鷶�F��1mJ=E/��(*{F:����BhJ�]�*z�+f�	���>�.?09�,��!��أ�;Eig����+��w�7�)����fh]��	p��AUBʰ����.C� �g��V2�?�N�:i��}ߤ����`6y�b��-���� h�^��&Q�鳡�����a���/ႝ�ݸw��zG��;�����KW�E�N�;+�k
x��R5�E�>�X�,�{��,��
$�l0O�N01BP�K;�犫Ҫ˛��/.P��aT����`�nI�$˭h`-�v��f�&2Y_�� �Mta
�8Ӄ��9n�p"��3�H��plG��-�C�sƻ*HaJ�> �tN'?B�)�!�N�_l 2�(FZi�(O�-oߦ�<�#t���@- �~r�e����J�Y_�'?K�i����Ր%+�6��� hd�g��+��:˙X����z�r�Ul`Ϊݮ�bG��Y^T�y��)sJ1bb�2���=�j���uZ���<.�Pz��O�Mx�>ub�GΗ��' E����)�C�@*y���|ūq#��v+�>D?B�<p�#��`�����Q++���u�5���t�g_�����W�~�gF.��B_�V��4�ڧ(*R��5���[X�	M�lN���A�NB�x��[V�k�m�i���(%�.�cJ%��=�p��&k�&��0���ԇ�
t���o4�J�FB6����or)^��@Q�y8W
��v�ڛP�������CR/Ъ��14m��@}\6�r�^Dbzװ��}X	{���0��90�ה}J�d^Q*
�<�����Z�4$�U�C�Tb,�a ���Z"�;��2�,����C��=^CB�`�uM���4>8���
�0Us)K��+sW��~RG�M�aN�&��c�}\��29ى���O���R�]xV���\�}���C�,Eak]#Ss	���w�΍���L�� G�=H���I�fL���1�"��i�LyR��V���0h�O����ȑE�9�f���w|�n�	'���i7�N��r�"�(�/c��E�
6:�ȍ2�7s�tڡ��a�.���w�'H%�l>p'�k0G���'�5���
o�S��E�a��)�3��,w:.-
qD)���2M�fˠX��:a�:��Ľ���N���G⥷�$��OxCM���z�e�)����71��xj��ؐ��͛LXā�ԿouxX�uֽ��ˍY:�#M��*Y3���b���[郄�qe�p�TWam� -,�
�Y3���W֮,P��Wt9uK����B�)�$�E3��v|$��Oi Df_�>���r��5���DԻd�����&��27@��"MZ����p����uì���͏��J-�ש#B�J��⹫��)�qG7�&�� ��B��@u����v���Po[��BCA^�doA��r�4%�Ӟ~��*b
'�U��k\��Ƈ�ih�����S�p�iy������g��G�3^�P� �^���\E��"�Ї0A����N ���͟N��2'<� �\7Ӿi�R��p�F� �г�g$�V�{|�+�f��Ԗ�kgoNn�>p��]i]x�q�?@<����A��-t:)m���*<ש���PY�����߁��0��0�[޹��]/p�7 �VP�|y-�(�/D�%k4��Y��rR�G./O���>J����?����Pm��T���� >ꋰ��-����#��;Ҩ(��	!C:W�f�j>b��љr�I�3�;5�d,ra��B��N9���MUԍ�b�l�?&������ܼ�t�ї������b���s	�X&��oP]�x�����-.K�o����0�O��%}E�+��f<Dm'�6�
:�L���|%
�U Ζ��2���#.�W��>��5�"�5�3V���,E$����]�~G�G�WQa.# j
��e�~vm�쳘��*M�|�k3�t�V�yؖ<Nmhr:�X�7<���D6#�	��w�K�@��m��R>�����Q�h�f7%���W��b%(�Ӡ�(F4l�E�R�����n8�a��ħ�x�.��,VW���*��,`�Xkk�m�G�J���06��>�j�E"e�h��SK�Iz6�� �d�u�d�?NE
�`=o�+���ZO��W�|����D�罩����G��mkV��K���ߖ����0�\ܢ^}d����rݵ��='�n�j�XT��$+t����2T��@v�L�#�@�̧�R�c��$ڂ,�N��,a�,���9c�m/��Y������Y�"��p^\�7N��Jn��2!�d����Iƥ��e�� ����$��#'W\�4�K�~~�Ò�i��W�j��e�/08~wU�'�c`�4w<&&�y�/���c'�!�5����G�tmE��Dpur��+������k���5y�h��o�����+x�"W0����م����"�+����a�d��"^��l�{��x��d��S�ҸG2C�}�U\*� ��e&y�����y
�岯b�1��"7���2���9xq�"��!�L���-P�`t�/Y�Q�nl�Dj����͓P��}��T���ߦ	�+��W�Jyd��ʄ*{ G�@|�����S�}�Ü���0R�؏OY4A����?�`��ӕ���#h-�r���'��ڬ O�;�i� Q��x=��~��A��t����c���y�Wƕ`�ŕD�=6aػdX�XNh}2N�}�qR*�T��im�Nx��/���<�
�6Ѻ���/Uҩ�7O?#�c��z6�;NeK!vb!�k�}�y�M�0;��H��fg�x��)��}��˖@�X1S�/�S8�L����� �K[�o��+p�I�T`��|�A��#�M�]�y��#5<�{�6�+�L���hEv�RCb1�-�v�Ǭ�nMZfs�?��O�xaQg]g�O��W�|��9j}��H��:2����3ҟ�y�M7��g�j�0 ���:�#E[�����_�5 ��ƺ���zy��lU���Ҽ����U���:L���9F�p�iX�c��8�j���  ��9m�N�p��KLh�4�]`���6p�F�wziw���H��dLE�z+��H���M��_�s?���>޶h���$(�i��o�\W�:�E�z���t,
�?�Ʀ�#%�8���w��8���t]u������f�G��h<���ж���F�/�vp!��5�����]�)T�@�|zc8��Z��Z��ؔ��V��G#T��4�2 ���:Q=�B�c4�Ir�!n�<��l3���:���J��i��z�������ޒ����H�.|�6I"<W�ǟ����fOA��|�+m�#if�a���,o٬�9S�#Z�y�a���h��؄�n|��=n�@!�)y�A�fQ �ǶQ�o����ь�4�Ր#crk���唠��h!2�lX|XF��?E�L�B��|;�-Lz���B��Ej'.��P>j2��˖9��m�M)�:MC�Ea	w��X2�(���ͥ��=ѼkS٫���Z����aC}�[3�
��QQ8���3�2lݍ;�v���\P[�z�I����8���k#6n������~Z���ǥƜU
��[����C�G������쾻�b�w���6�k����,ZZ��b���qN;i�4p�?`%»U�ll����f0;>�hg��Ew�v�.�_�?���>G\��+M�+؛���y�h}�_lМ5�eO� �Ǯ���޵�/!?�X+�k����$��b�p~;�dc��T�ykm6�@�������K�!PN���F�Gw[��"2���+�p�e�&�+Ѳm!ڀ��n�#�Rq@�b��@4M�}�B��t�TrԷ���5��N#s�,o�d\:���u�#�-s𭙕l��a�s�k�?0������݇g�L���Y&#ů}�좋 2��C27���Џ�+މ$?�FMw�l��V����|����߽W�!���g�R�w�,_9f�|��m��LM�M�hۭ��L��)Ʋք���1�	�����Ye������@�3�B:TP�Z=�f����/�<՚`t��6�g/N����:�ԓ�%��	Vz�fD�ag���S����[�I�����oR��3L���AP?c����@[ο�C�w-���''�BZ�6Q�`���s�4րKl[�x�as>.f���P���\����^�A�A۩�ܨ ���c8fE�c2�m_�HV觥q\:!�9���h�Y�#\�.e_HY6���ӱ��w�64�����"�J3��]�V��gosk�?2��1/���� L��`+C,�
 r��u�4y��]��2)��۶L��J�����>�8`i���,\j	�GJ6��Y</U◡Q��ţR�����׀~���2�_G�|E�D�tÍ����t;=ҕ�AR��3c��ݝ��)w�ذ�|v%��"N�h�p�P���ExQ�7's��-���{�Cj��łvk��y��/�c~*��7�|�������jcLO*��P0, ^���a�&s��[���Yl`G�}�
Y��{�@�U^����(�b�=�Ϛ��&gu�*��~'�k�՗��O��.�����מ�f�z���2ĉ#�[��1�kL�@1潝*2��r�����u&0��'�(�IR��@E�LD���z��d�c.����0`�ٸ�g���{=�����2��'�h��a%���W�� �n`*�32P�ҝ��d����qF0��%꽫���4�ܰ�e?� ��q]� n��|P�1/}��ӡ©Z%֯�A�� ���i�Ĥ��1 ��8���w��h4�	��Ɔ��ӆp,j�&�5�Bz�<#��$3�Z<�
c�6<t��G�� ���Y�E�#,�S�jZ���j�T٨�a��!� �Z?x�j:#��PM�kY�\c��Ie�/��_�����e=6Ud��"xH-k�ڜb��ç�Gή��q�<�-'���$��������0�?����1��"/j�A����3C|B��:�����@5��u?G�cj�S��nB�l�����)�����āw��.	�]!�U�N�SH�k�e�e����bSԑ�Sf���Xg��k�z5�v�2���#!>���b͍����`=�l��M2	�9b�*��,c�����E<������{�i��!�a]��=ch��R�!�CY6Ot��_�E)�1�0��0��Aa�,����|�	�އ�z\��m��-͉���E�7�4�{-}W�O_��kR�p���G��8� ̮�|4/Ugd��'�e����l/Y��*Ccۦ��I����e��i�?b�3�}�u���e��cfr���ݠ��/�0�"W՛ }d�^�pa���\��J?�[���8 ���A�d�Py�{(z��1?��զ�Ǻ�া��ToҹC�H�p�5��Vt[;��x��6ƨ	��{��N)%�7���!���d]� dk�9��W�nHyGC�������6��Q#��Z �g9�T�ʜ�V��W�HZ��\�`���<��ApW��9L<_����Ү��w��~���/�3�ᐷ�A��5A�x�`�m�ՙjQ8��#�tHb�>c�p.&M���%Z�l���������O���	��XM�1�G���|�M$�B�>��Q���{�w���FR�?� �WDoç��)-3Q�ϣ�$�ɢ��k�p�pFs�W���Ú@Ԭ+7����$�W������M jK*'���R��όz�S�4�0�ZF/vjB��2��Y�Q��X�0�N ύ�>�lᑐ�$�NB����C �A�,v�ˆ|sjWB��vT�\��I�v4z���ix�X_ge0%Rt��4U���9^�$߄{�s}�)��~�ߜ0��(��8�Ң��o�x�z ��Y@x�&4]�EO~��V>c���p.۶��'�5-6���ϵ��׾ 	�1�����א�J	Q��N,S�ik��ׂ�H��@:v�!���K9��� S�w�i����ȶ��"�>�Kk��ۏ�HF�ћK��L]#*���e|�E*�#�ָ9cG�?t,��F��6�!#L�BX,YT��2<�gy�#EV��85_�Qu�G��rTtܮ|CF���6E�;MM�⪣�����_����f9��ۉ���1Zm7�y]���x��z��rb�G'������)���@_#����r�Ǵwx��wR����D����.��*�����W҂�
�.���)�+2-�7�&�w��/By$_G%RYDΥ��� ����]N�H�V���n��=R'*2lF�tڕܔr+����6�Uq��j�!��v(�Ã��1�����4��>c�e�GJZ=����"�����tβ�b���PC��~"�֝�T�x�����i(C�y}�Y��w~RK�'[�`z��EG�)^ ]�A��x�����"�&�%�#�m�5��\];:�=�0�B���?��7��3C�-��5�{A��䷔I4��NN���U�p�Fߟ�N�Մ㈶����������ҭ�_�^�(E\^�d��Gj�U��Z�H$\+��:Z�s��m]ƥ�Lk�b���ԩ�,�/a��]0�,�nmh'{�sJ����Wa�d4�j��J:Ʈ�{�a��x}kn6������2
#ڑ<�,���Ѥv��ze`$t�s	��9	E��o�!�-�x�8��M�r�	8�q�9�����*[�<����� ���-���SF�Pb4;��(��F�c��	�LM!`�|��N��ؠC9BW����]c��M�?���n1r!�O�F��P�k��_���h�ޡ�:��rM�0�)`��� �f
5���ϥ��@���t��#������7�-<�����"~��� ���m�{4�X�0a���Q�zH��fuԏd?�y;JF�wx�����_#����@�9j	�M������ˣ�#�F 2+��x����a����0t�Ƽ�ǘ*�����QI�v�P3�t)S��)OHc�KS+�p?
��K`�<��\4>U�Q�_����ZC�����
��O�
��'�йp{/u�壘U���&c�S�<����@��{�ρ�x2��f܉U��K����P�B��g��M8�s��d�ѽ."e%�&ȷ!��XR��E,[f�܆�)Q�G�\���,���(�N��l�\0��	�ĉ��<o�0�w��`��.���J��*ub�ihV�P��"�T���;��Y�K��� I�Ι�C�H\Ŝ&�^qN|�)�C� ��|�F�v��B�A|_����j΢tF�YB@F8)`0n�)H��)7V��^L�`�e5v�DX#�X�n��5ÄąD�r��]���{Cm�ͼ_�t���o�"�A}>���\3�:�w�c��-\���Vs��Gy�����[Q�BŹ��J�a�����h��(o�"+P��,%5��8�@V�|C�������Q�����ư>��%���d0���Eo>�.�:lZ�iQ+k�Z����M�hn̼KX�N�P����"�36J���g����Uo{yˈq�hx��fQW��a"�F9}4���q��͔w�A�Q_�� ,����A�ꈘ�5e�����@@v�>O%k!5ql8�f�����S%����]�X��5�z7���˫hqti�2݂�9��{��c�������|�O��Ø����P+C�Ő��I��͂/�n1��ko0���'v!R���(��"�Է�/(zO���d�lu�}���9�E�2T��]����P��|�@
��sGHw�.�ƧOU��P!2mD�� �����u4�4x.I��K�	�T�w���/�BEc�E�2v�8	���T�Q"`\ ��Ν�єt�9[�XD��w�/�x��lHk�W�'yb#u��eY���ZI6�u�U�e�UѢ�Ш��_m*ss��	�ü� ���H��R�f �J�|) ~�C������^_�i�C(5I!zV��A��>�`:�h =����R���+�9y�8gꐙ��>ʧ��a�#��`4�̆4���wy5�y��nf�	�B��Ғ�I����c"܁k?�\��M�Ys����F`��+����3�Kİ�/��'�bq�0�;��"�'�����	p��8�U��[�	_2�<p��A;t��m��8�4��J[��#�k�=ݾ1�g@�Ԩ���FJ�gD�䑈���ע�z����2P��Y�@��|[`�)���d(̀��1ʴ	��>��.�A����|,�T�#�~���G9/���^���"���\�f�%����F����;�4��#�74�%�#T�������K�X
yɳ��@d[��!hI��d0�`k�X�r�ST��W]�J;7_冨�X���-�	�F?�F�����3��\�Mp�ƀ��v��
�����#.�£x�:�@y(�V�#|҇�b�fj���'	�g�!nCܶ�2z�&R1��>2,!���η���mSt�"pԯ�%q�Ҋ�P�84c
�ƅ`�#���o�WSp�*s�%e�{�0��̸g��,l��j���D���U�I�A9�6�^�ڄ����D�]8nv4���Q���.2�y.�G �����U���{����J�(���a�cn����r��If�Tl�j�6�5��y��*��>vC}K�5}���'�����.x�7͐)��<|I=d?&x$�U�f�!h��c���at	�X��Z
�}�)u��$3��W>�,r�J|��mk��{TBx�S���Cm��d�)AN��v�p����/R c`M�>:�4�W�Hx*�M��q��Ʈ����U�&�/�0Z��3,������s�u���'c �F�ӽ��-6u@��w�"��C���B&�׵m�Mw����?�i[,���U�l�dAj�` b)�"�������� ��]�A9��]v��/�������S�}����2���(sC���|�� ��L�*2�F�i5Q�R��O���gtF�q��4��)��W�e>Sl=���L�`�����묨�*&�=E��!�[ެQ��+:l�|�>��\�$4DE�x^�9����'�x]��2�o}�w,�},����7��.�.-�	�c�^�^;�ወ����|r?���$���x�T\�aM9���a�0�4�>E#�}�8�O�K\���nZ��v2��Q�l"(F�G�8EB���B����gn8@q�m��u�d�#���6*���!�]��I3�ZuE(�{�7ms��ɽ�ؒ�2�s�[�'�N���Uid�-���bмW���2.�H��]�7�}��+#-l�^�Ʌ ���6��dq��h\k����{�GR�O�hr�)w̿�.�~��a��� ���ꠃW��)��Ц*	#��`��a68�!��������h9taLd�NW�ԗ�uQ�%�o{q�S��0jb+%?<�U�(�$�%!��4L�ӝ�N.���g5��5� e��]�V��j��y�|�T��i)[[���TVn)����ڹgX�x�o�Ʀ�`V]%@��a���9�;P���r�m��*Й�Z�tÅ-o�k���n�,��L$L�9w�m����G��V��A�v����+}Z�ٞ���|k����dU
�zw���30���L��9!�BIZ?�!E��gc��H�l�N��|����}U��ق��G�$��{0�,^6�_�7�r^\��kf0�	����6¿+�S�c���
z���l�\\xN7hpy���?#ܬ�������hO��I\����	��6�N�E9�<�6z�@�Ry��l�]~���!3�q��
̐��o�sd� �HU�|ryw���� y~�{���oqFz�|o�z���s-P�w0���k�j��T�l-딢�M>4Bȫ�Oߧ
�T�v����uKS�$,�����V�6�2E�k{�7H����WC��c=��!�!8�eZ���%��x�E>^�>(3%�]�*�餜��rV}�i�C5��R���� Ϥ���,�s����:��J*GX��>�U{Gi0⦸��Ǭ(�1}vq�S�*�!��Md0T�'	���F��C�d�V�4�R��Ƃ�^�5xWv�_��[50��H,Ζ������f��٪�w�Di�8�Dp��3ɋ.���D�w���mfCu�:�G��4��7%G�P���lː����O�k!�=�q��T%�P���zgy?=*܍�e��W�2Y<*��'�2��Bh���b�#�w��)�А@�����0��M���̔[{
�ڭ�jI�L�mᬯԷ��y�Su�q���3������.��U��3$�6/���(S=��ky򐽝��ة���1UH�:��T�,;̆�V���; ˔*�vM��-��D�qT�r���'R��Ɂ�z��3l�R�?��n��QA���{,���I�f�l{�Lb.vh���Fҥ
�+<�X�pu�ܢ|A��'vO��l���7���zX�|yg���]2�i�\�O�?Յ�~:H�C>��k���ף�p����!�Ag9~j��z�a��e �	%��V�+Ύ��^��%įq[� ���x����+��B��������ow��Z�]�Q���H�# x��馬B7 i\.����Kz�5�p�@΃�ŏ0��g�7�Y�6��.�6�鯐����"[��M~�K���z�]�R�`���B߹	�Y`ov���✤޽�W�ז�n�m�hX��V���)��s l$�&���-uDc�ǀ������W4�Y�תz���k�>����ЍH;y|u�F��$v�L�)�ؘ?/Qq[��{_���$--���]��v��u��e�)d�դPH�9:�ɩ��L$���=
�{��C�I#q��d��Ϊ�����E�_w�
4����`�q��`�A�������P����T�w��>>fz�j��7�:��B�(V�*U�C-k��<��(��Q~U����}.'}�.4���mF���y�5d"
B�7����!V��l?�;���-�Ж<�L ��txd�v |�:�kC0\YQܿ8N��(o4K���㨺+B	���՝�j��aAr�����i��_��E6�
�̤=<[මH��qN���٭T ��nwu�|�������q]/�l�z!s��mhO�"y��V�n�)P^��c	
�����ɊO[���VrI��-��z��*����wI��&�+�+
�}��I�'�v�L;����lVzw�Kp#a�g^2�}LQ���&��b�'�qb���t�,̲��: ���U��A�����7��T��*��i�pnǒ������L��=�+|�N�Hsߔ-]���3�<��h�����@hn���;���ِٝT�����SE$�k��B���3�DD��"�~%<>��f@�q��XN��!s9�(�-~�ө���ߝ���1�>;k>�ʱ�t�A��J���ch�Q�)�}�0�+)XY��7�ld��J�;��2� �1�%�ķ:H��
�ڈ���F}�f�k�[D������4�(+��x�Ch�+�d�=z���ŉ����ȑ�J��\r��T1��/�ez��0_+4;���'��δ�D������%��&{_m�hR��, �v�"%���	�=����� ��o�3��5ѩ
Ddg��jS�9P�
ң��ή��J�����.%hv�7�o�dR{��"%�{[��Gʋk���8�S���1\�����|xԴ	�-u7$h�5�Nb�X��1X��e-`��7m��G��u�A"��ϒu+����I���$�ċ0� v�C�ۀ�>u���?�������"�C"�¡�*��徔�oV��j�/��!�q�5�����	���M_��H�O�t��{���m��y�)ss=6'qB��5�=�eP ������@�#^��2A��GZ�M3�K�����Z!*��9tp�D��Y*��K�`�?N�'�+�iz��V�qz�B,�rGI_n����.x�oS����ms�ai<" ��ʄd����Z
)��kŨ�2�io�S�i�zr�#L>	�y�jל����8#~;�D�X	��Fާ�ٞ
m���+������d�'�'aS5s$�i�K�\ʎ(����Ps��8��,���Q	vz�G�ُ�.4Kc��@�ڛm'�O�O���w]a��PXaZ���n���`�@��П�>�������~E���h�7�	��!V{A2��,-88�ȴB�
�]�
�t��=r��d���$8��+Y��.�s]Qv���֎���y�����(k!ᵈn�� ���Q��!5zfI�8�;3�1K9
���.(��ĝ�O�c5W�z�BM4d�[��^פ�V�~��� ���پy~�7y��h�9zb�OM��:�q���0r �(D{��̑�F̿�L�f��-U���Z`%9�WK�*u ��H��|�*+E�.�����N��[����"�Fry�3�8����>*IW���^�zu�FҴcl�Mz���_+$�S(��L�%�=ĭ�]��0�u��#�Y��D�Y=��U,�%�Q����R�I�u=�6���]?��`�t	���d�@��
<q��� Ҹ��x���˵LA�����B���h����Bo��ᨱ�p%���R&��q�O��#2�Q�p��N�&q���[C+�`�k{��m�Hc��B!-��~���ײ�*��vF�P��iA�ƢJ��I32]���&N:xW�u�}�-����am6U�K?�؍۲W���ɤP2Ǟo[�@�,.�3fX06����)}t��j���Dn\Nn�@�\���șv���R�g¯�F�/�QB�/����x�,sO�	t�f�7�N>��P?u. �vs��q���:�t�>��� �L��A�-�1���n�k�u��]�����K�rI�w�L��R��K�&ܖ>W�α�V*�/u��!ˌ��Z��7Ѯ�
�x�$G}�t��L3��]*T����+��ݺlHؐ�?W��\�F7��{���q��=g���@ �?��V<lJ�$<�q2.Ԟ��Ž+	�������үe�DM�F�"ndM����Xtph*&�I�]���'��0{���vH�]h�ٕC������w`��r��%Ϧ�(^�H���˭�\M�V`][��Fr�B�C%j�3T*v�<d��J��L�o��<��X�Q�5�ȁ�"���;$싍�����8�{M(a㺋nܻ�m��h�yо��ȅ��.~����Rr��y�i(|Ǽׅ�uA}�B�-x���F��3��-�k���[<Ϯ���ȲA>�0-��zZ,���Km
@C���Aҿ�9�8��2��r&G!64p���,���.��� 8�墏@��~5�u��әg�B�����)t��`���
E�3B�\6�#��sa
u�f'�^�и�`M�{���s?NP]����>���Ky�����s��{"�b���s�=���I�����D@L�d�t��	ǘG�?��G�=�Y��6��0��E��u�
�PErwK�\x��F�!�����`���O<�B�J���Ŏ�J�ar�v����4
��aC�Y����_�v�2ޥ1��Mk�!y������P
�ൈf-"�W��+���0nc���0,o#�f<�����B��AG1rm���7.f�^�1H��7����']��`6���d��S�u������!�
@�����L�٤w�#�5��F�v�"HJ-�*(���z�(E	}Ot`W�%9i�T��Hp����6�Q���|8���~�!�^\�=��y��Nm�Cʖ߼~�1&%9�������,3V�tЮbLf�7�]���BëjԷY9�4�^��"T�F����/���������H��u� r��)�5(��$���o��)���Vm88�:vR�v&�z���fv����j��o����i'?]l����o�IO{IeF�(Z$)H�(���j�b�,��0̎_TO�.�xa��T�����4�6�=�Mmڝ ۅ���awܙ�N�ϳݘ�afR�%�6%ҡ����"�Z7G ����(�A��-�^;I����H3�������L�P�����w����>gV�el�P�Q�?�"}�}՝R��C��.Q35�>�[e�!{E�d����7^ȟ���.B�x���oM���Ag�P)f��FѿX~֡���N��I�������B�_�k�Oyf��A��#_\Bg���P1����%R�"�p�f�0��̤��'���^9s�?RUc�031����p>�Oh�m�#�6D�j��8 r�����o@��A1�'���4�NSU�w2������N�	z�K��kd�MR��F��Ba?��Z��x瑖^�-����{���%{�ȉ`قa=�	k���4PW�nq�|ó|��ą����&�qzG:gY{��J��7v-�V��T�5��X+�^�ߚI�� 
q��*/�ʗ��z�Q}�����۹�$r�f���_L�|t�wh[�S x�Yb�gj��s��9�X�L�r�zK�s��?����.0ji�e��E�ee)�����q`�Ʈ�ϰ.�,�8YaKA�}���� #Jx�U"���:b��<`�{'c'�}蝍����<��'��Y�p����Vo3��=oN�����4w�'_噘�I\�;�
��'�J�w�"�Oe�����NHU�z0"yh��6Ӵ�)F��mA�`�V��xB���5��N�xe�"�����
jiޛ����)�o=�L���R�h�)9����������5�[���p��{7�<�<s�X璶��!�b���<��J��w���	���/�Q!<���75%����iY��!��z��
/#4FE�z/ɴ���E�ṰO�k8~N������V��
[\�{�[������V�ni49��8����T;)�S���⸗� �K�I @EQ���[N��}�!faG��'�1DpT���n��Y	�g��@����Yk�(��@���<�xbc���b����տ:Xsp^Ow�K�Ҥ��C��F���.?א;&�%Z.�4F�Zu�a��j������m��iZ�Q��
X�pzD�nt��xŶe�4������bBL�r2'�F�7��a�а~���)5*�u-`�⥊��2�͘ת-^��b�ڣŐ�jp�P��;�\�j&^���}����ݞ�]�E��#@8�*����2�U㕱�� 5�II1e��a^���"�u��@�4�E��%�0H�vX�c�\Ob�_P���R����}��;��2Ȃ ���/R!��7@B�'޿w�a�ݵ^L�x�J��.P�x���������1R����\�	�]dS�*�����.�*O���aH08�Ch��n
�^�����p�H���U	 +E�TI�4R��Ā<��6���pacv!������u�7���V�0�"J>Z�K��������YX�}�1>p[ ����a%��k:�N��ɓB΍1H�U^��'��/C�j�n�GGb�S�G��!N�<� ϵ�mܣ}5�_�F�	���j���Y�`!��%0���$�|�\���$oZ��ڲĎ.)��9U�d)���e�W�]�.6
7n>� ���i՛�xF��~�N�u21q�	��d�OO=��㰅7%."�YVs5j�l��x��;4Y;��������R�)��ŀ�Bϑ����4����]�Aw+�rK�i�RH�=���]�NI}V�ܔkFɝQ�ܮP�y��"KD����5�擢:�L>ʶ���W��@���n�E~0d�0���=���3����]��\w!X秿��|��:z9	2w^Q��'�g����nb`�i5�uA��%��Gs��B�nw�þ�e���}�P���4�+�ћC:���hE�Ix��*�mؓ0ʑI���IV�#�B�a�π	������n �4�E}z����%���?����f���M�i�nd�-I7�
h�h�冷�*[�H������Aez �Ɨڍc���+��2FcϢ��A^yU�� �1܌�U�z�.�����zH���� PpV�I��xq���YD_�w�8�h������,��C�ó]H�]��w���$�(Dw��D+����Y�
���PJ.�s����|'�J��\A�q���$�Jۀ�>EP�������}�<'/�~ܽ�q*��`0��"�lKzu��Q��ɹ�J�mmc���}H�33^p�Zy>7/��K��d.������
�UR�a�'4�T$+bPgr��6��j�;��s�N"�⇪�~��(ٌ�'̡��Vw.뾵�x�SyԾ�:�OD�|$g��s�^B�!�kHsY���0�����HȞ�-Xj�R�`�d4��K��-�_ 3Aj�+\j.t]I̶�a|7������t+i�#f<�wԗk�꾛�:&��|��Is��������冝�~�,BĦ�Ɔg_�!^��?�]��T��7p�����6�Nk�ދm�a{�͌�ڱzK�K^�P��֏��C�O��⍻.
�Q=��|f�����P%��x_���K�Oj~H*W�l��ԱQ��ǽ���$�؄����Z�:J�v���:�8<�8$);u�2��������7cU衻��(�ܥ�`�a��V��D�"D,j7M�E�w����ϫO���8���t�+#>�]c�JɈ*+�I1�_�jGIKt�5�$�n�����3Xq��gKK#�<,^��u��!{���Z�5��Oz��5MK�R����_�3��cu4�d~���tp{����	VO`�K����k����e;�!�_Թ���@};��&�A� ��:Cs*�r����i�][���V-�~}��}<O˫�ѧ�G'5"��j|	�cU��';A����H߶]x�����k��n��|]L1OP�	8ٔo��"�Ӷ|:~+z'�y�ǯ�}B=Ix���E�1�b`�bA�s�ug����/l$��)���g�(��R �E��%�{��g-�������ֲ�2���]�c�gUE�x�A��'�MT�T�i*���Z���SIZ�6��ı�
�{([�bR.���q��c�$��-Z.p2St�.�%Gg
�!�)��χ9p;U��x
��B����gf�#w#���e� M�*ܥ���G��v&�0�~S���yR� 1c��o#	l?��eG
�>�)n�0��;3L�_j?��Q��I��i�M)Z�Z�҅u�6����[L�^�;�g�`�ɴG�L�X��3�q"�(�@��y@9�'*��Y��;�+��' C��(>H�L�G�����5���kL ���a�Y@�v����C7�Y��dQ+�1 ګԆ[/v,tϛ��M鄡~����H4n�՗\XL@%���fy�E�WD��eY�44���cM�]�e!�4K 4`M�������9��pa�-�����4�IR4i���䋤��;P�yg}���QB�@6�0���
��HcG���f�J�����_(�!�b}9����&؃�w�n]�X���[�5�z8��XU�X`a1�Φ ��oT��3�a�L���ǉ�+����cϛ�{�]�Dc�r5�EZ_��D��wv���9�hq��؋����G&T���Y����v�	�Lf�Zq~�.�Y	�*넦��6��a���/=���p����i`��5h�"O�A���#54ؑ�&i�7�0P��`��n��J��_�|�"�b]�"rԺ��3|��RB��p��b����1�*�|T,�d@��`��y�0��i�l���6`�䏏r��BK�6q�H���!�L�g4��BZ���(�1��0}%� �^&�b��+;���v�t��Ʒ�N-�!�ъ�N�(��hH�������H����G#�: �O�Aj�fybdz�E��.�
�8��a+A?�����(pi�;(�HgD�Z���S��)�踋>:���/E��`�0V�Öna���(}Ҏo�=v�
i���f�����x��	蟄"��.շ�W�_����m�F �߻�HԪ�˫uT䥲=*�VM
ऋ`,J��
uApX�Ne�$EnG�{q�� )�O�<���9��4#��~���`qk���F�	���|� ����H�A}D��f������]�T�:wV+����G̨����H<��4���DKM���9n���/�s&��2���U}��4��(
/�"�t�Iv ]ւy���bk��^>]"��J�_�-���至zo�1�x�G����Lꎺ�.��π@���؀�{�&�e3��˸�M{�+�����S�A�!�T:�mxpVE���C��j��f���h	\�#���Qf h�'f��B&�RpOn��0�B��H�]�G��Akv�2A��M����6���p��t/�2�?a�}
�<C���ԟ�/S�y������8ϪS0���<�^�Zk�M��	��]�1���^L�7�a�Ǒof!q�>_����1�@ef*�����J�"t�����gO6� �ܛږ����=��`�q�	X � ���cV/���ZI#��Wfҹ��Pη]Tj#_���Ƀ���ԅc��Ӛ���cb������`J.0!ڞ�l�m���W�Z&�����%پD��bS
�'�1f�/�U�@��ɐ��̀�Dx��&6L�o�_;ͤ���2
�q��T1������f:��
�� �&�K͋��<���xX��X�ӵ`	�j��6�¬��2`�4wp�OLQI�z��vՎ�8��@��X�_Pl�Y0�Y:�=�3.�q�9�^�����/�{��eUm��-HSV�!�C�����o��N�v�]	[_�_] ^u�Zk��@f��q�����e�,%���R@�)��}��,��|�BƓ���![�!�&r�)=��1�|]Pvvnx.����߼����OAФ�F]�Re���W��'�D���Ux��M_kK6�� ��i	%�V�8w�/�E�<��Jax�}4�b~��������a��x3,�!�ѼMx5\�4��=o���E@���i;X��ۉp��]��1>$F�5� ��ZX��qu]�8�۞o	��Iw�w����w�Ű�ޮl���l�����F��T�#ok�h�����1]�������͢ss�;�^��m���������pf�:�A+u���Ӟ��J��.k�Y49���<�4��4�j��6E�C�8�;69���"��25�������h�Bmq��z�',NkƶШ�A��=�������PC�n�E���g��)�x����_��B*�L���_]ʫT���(_ 2&{]�8���3�0%8p[n���n
}5l���qi�](u�T�@e�'_�
g^�Z�ϚoX��WNk+��m"w\��8P��LF�	��:<Uv� FC�+PW<�J��~~>Ɛ�K������_�9�H��hU�DO���$��68�yq�]YE:a~UQm��cR���3z�/�VYS�K����6�Kfj#V NhA�t03x�Z�0��^/��������[�g�Ø6��L��u�3�(�j��l����,X ?Y��y��)��'�A��E m�Oo�x��_��Y��%����	��l8�j�I=�9u'���z���k��+O��q�?���U���)ڝ+w~�ujQ�V�a쉀E��H�._+���Ǟ�̸5�/O>f�����=�F6m2L?�̑�9����%�� 9$ c�7���u��}0So���m�X�>�#4�hT]1��?�=�����-

�{��#uw�?

�`�ֳ{��F(��ln�g�YYw��D�E� �<�Jx�YR1��ڰe R���^�e��8�#X; �����xӔ��M�.�8�k<�q���[����4Zپ�=(ROp#��{��{7�3m�f����m5�ϑ�Яڞ'��ZRlOa��G��e����e��o�*F��/�K@2����^�.���[��1�}�G�c'02Z���RnY[�pE^�/��ҡ%8�+���tt�t����Fmֳ}S/ƍ����mJn���H����
��EC~�޹�#�Zv��������!D�R�DI�7��*��"����X;8J��G�@���SR�Mr䍷0��$V�xx^�)�쁆�l��A�w���"c�y�� Xk)�tKF�թ|q ��:�q�����«I%��t�AO*���Ħ������z� .�F���	X�d�#�� 2�eA���cz��wgv��
I����`-s��9�'�0�]I�Y~֘Ǖ%H��Ӱ���e���l�4���]ן�J[���ր����s#$-Y��c�5��tK]vPsS�"d�@l���oɛ�?Cf	��[�+kE���,��	L2ok��-O�EڄGGGs�C����ƵpQ(��[����/�8�z��F@�qi�d�]���7�a�o,�z�7	>�o��Vwm�2�[���&�\�z��v�*��y�液񳘖r���������4����V�;�SAr��c��6�,��*��x�Xg2�q�t,�H#�d�샍���JN�'�kQ�J�+�D
�t�c���D8�j��>��ߞ��������A��ƃ��-��������v ���h\<L ��q�E,!�����I��p��1ճQVӸ�L�x�f>�ƃ���>������>S�A.T%�2 H�VM	�ur��&\+�]S��
Br�
��\:��'�fo�u�O��nMq�t%���~s�4�l�YCt*#����J{Y��]Zk�E�,A�Z?�<���,y�4�?�x�HQ�@٨K(yĬH����H��자U��3����Î�6��h3��z��.�HIIn���cwY�]"W&�Ii����.%���`�ZqW� !G�R�r>0��J���(2��DV���Յf�O����Jb;�3��s/I�5eZ��KP$n��BӨi�;{q&���T��l�Dˑ�;��!�kK����,܊�,.�_�I����e���k�B�!0Xm��%��1#��z9cC��t�0����󤂙7XEZD+/����*R�I͜aSu���:�'���¢ui����6�>"�i�yq`�L��FD���.����]��k���\4yݛ~{|��$5hH��6������d��N�@�� �{��(���h���3�_0�������K+���6���ɻ�S�i��j�kv��+��9�i0���؜���̛�pp�b�f��!�~�4/�9ԟ%7-�depJ��JN-�E���x�;j�-�}J��}x�hi�?���_�����!��j��1�4�2@޷��U��&��'�������RV����"�%�9���n�����:l쨷)������;�ĢY{��Rf����c���5����Y�cN��dƘ������J�ll xJ�ݯ����e8̣�>�F����A�}�ν���y�1qF��ӱ�����,�I��Rt0_��S���P�D$u�ΝE�vt�/�k]�=��V�Ҏ�O��e=�)O�+���J�A�x���S��Ԭ0��ű�a����z�n��v~a�OaHvU%gD/������q>O�
=��&1-���� σgj�mЮ�Q&?����&&_:	{R�+�j�]l��ʗC�_<Y9����`3�BV��{�� ��_��N�;5�j�����Z[/]y���5�S!?a3ñ�O�¡���!��]�J�<M��7>��A��! ?zԛ68Q�Z�}����*ep"*��?�#��Q�ͅ#��8�\���#WJ���N�.Z8^ͭNE��i)?�M��.)("���S2��$瀃8i�&<�Ņ�f������@I��� a?3@=�����~�:))K��;��5��ǘ��{�6��� �AFd6���T0�.37��R��Gpcݘ ��=����Y��t��f�V�d't���P����>l1�M�s�_�:nF ��3׋�������n�nd>���қRa.�<��큘���h��ˍc�ne�q	fM��Wۖg
���z�} �0�[%�l��`����i�Lu��=A��$�b������֪�se*$ ����N���w��ƃ*�a)1� �N<�X��Ux��w��d��Z}����X\�4s-��܁�U�jܹ�H��$F7B���?������0C��k�M+Iq,
�s��t}�@�Z4�,�{-��V.ܘFa=d���O����x��}ם_뱝@�ڹ��4���[~&�h�������g~��k�|���m��{ �2�v-`�21�ȁ����_�NtxQVL�D,(���17�k� 1"��f�k9� Х��X���:�ͣ��(Ҟ�VBb�'A(F�E/[^���Q�� u��#�d���o����=����T�%��VWw-T	ou@�+2G,�"(�1�|���n����d0\u*1�GYj�Q}�l�KHQ*O*��(m��y�7�0>%���ȩ0��f���WL?M*69�lAF/�<�vD��u�e����*3�z��m�}ϴ����OL��t�8����
�U�v�e��� �Ή�&���9�ƌ\��Ҏ-͎jY)�?��V�%��#�����e
@��[�4�����x�ↆ����ڛ�B��bR����h�@}Q�;�,��eUS� é�Ŵ`�_C�~���qX=E\U[-N�>w��{�����*gi��Plo�Y9�%k�%�����-�Ξ:K������"`�4����io�Q�\�)idk�V:���Ђ���ٴY	o���md�����l5:$x�ӹ�1j(�����R�o��9�&�^�>[F��%������v�ܱO���S���|����S��[�Q$M{^�,{��q�#�4ԫ[5�3��f�m�śa6l������+o^�	�˲uݍyG��+���$9g%U�}�I�C�0l����z�d�=k�N��fi颲�g������f�&��B�!�rx{�?��,V���C,��Y�"ݼ�kS���ˆ%��M<�}�p���E�:�J�;�*6>�)�`Q�����g~=�yџ<�wzke��ec1�|p�����
K�q38hQ���Ď��鎌"n1��(`%)y3c4W?�d֮~���9��#�3Z\f̔R9/"������@���lEbq4�Jb���7����qv$َS������uP˾Ԋ�{���⭅>z;�3 ;B'����]x^ͼ�"��8n��d�=�����	ԛ~��p�� 4^�S��fZ̀���i��z}�9+��^9tE��P����8��Ԭ_d�j^<�b��DS�F�Sn�A�4k䓎: U��?��x�u����<��	�rCP?>Zu+u�;����۫mA�Fq)���>`^� "��9%"��O4c߻a�[��r�ׇ̗c&��t�y�J$Ro��;$�ۢ1u�P�^�(4���.@�%E��Pp�x���m��-y����@_T#��ՂoZ��HF�����p�C�?E�\v�NҨ��:kg_��.�y��^ԤB�!B��cbm�'������p� :+t��\����f�� "�Sۅ�����~�q18���wƀ�Ӷ1��$���-��G�>�d��vIpc�R��=N�7�������/���LRO�r[�>f�L����FB(9Nft�YU�c�Z�Y7[�N������}�Z5�����y�0JN%���	/�ʸ<:Y������w��ȓ��'�p�#�/���C$Ǖ.cD�<EA!�e�o�-Fls�ڹ�$p�6S�`�TOX����j2pIN�uѰ�b�#62B^��7�e!�������	?��*�J�� g��.��^��_��¸������h�Vt���o�Э���j�d��/��BoW�?�[��{X�2��Pp#�RCC�b�[��Q��U�Ʉbz[;���&vh���X��m(A��9��4�.Y�&���7�r w�=��$���cV�lܹ{��$⁘�[8�7�?R��4<��yf�o��\�9Vm[ku�ZGg\X��L�,J�&Y9�L�z?�*���x���g4Xίԑ��B�#�Ykd�/p�[}�k���:�LK��0k�/ ��A��Z���U(�e��$���%-�+{�E���5x-�<$s���A�o�8&�+�>�]��_���(�M*M�7CUV�0��?^pp�����s��/U*��M����R�3�N�c���r���3�=c���B-�n����}��P��h2-&#�V���i_�fsBM�h�>`I#L��Az6X:����_�Z`�C�������N�8͉U����R��ٔB�_EbƲ��Z�ƙ�]v��q��G�lc%Dx�W`�+D�1 V�z������]��ZU���{\$"���)3/���Fbs�,��0C�%RQ�l}4�lrQ��ڳ޾��%<�<��Sy���W�<f��#Q�*	��c�`�
�D�G1ڰ�r�0���ߤìZ��jI��3y��[*	�j�ڊ�#�k����li4& �uf=݈z��<<�r9v��-1�_*+}�Z1�~�`t�����Rg�3�Hb^쌨#�)��]V��Z�ß@��W
$Ź-����3��h��ʿ{ظ�uv��uG�!�)p�<��\A�x`M���u{�PqVy���?��MfX����o���B�]},0iꃛ>����$6Y����z",O>2W����W�'�_�2��:;��VW?�9U;��wWw��@tw(h��`�iF�82��SȐ$��5b�|X�T����[�]�Ơ�T�L���D�3��A<�l������%�2��V�2#F^�X�{�b�B���|�x5t�����[3" �\�	̜C��q�I�	����<(g���s]�HB]�S��1�+��gInN���fu�Y0���V���&�W�f�� q �f�T�!�M���m"�y��B���ˈ�T��/��4��v��|�xw����R%jz�
gq��翾[f�`�P���t�H��j��6���k9~�o{ɸ@��$2}�fؒp�{R��>^��40�r#"8ò�?�c���GZhN31���h�&��A�ݢ���n��h>���\��W�e/9F}"��&t^�uzў����3��]��zc����M�����-�*���K������!�����yhN�wt�C,�x�9|���4����`�؝��_M4�y�54��.�Nm~Iӷ�-m�[�+�'��@MYpԫ��_�����*5�<���'��>zq����S���+�����L���e0	�x&��k������g�u3iky�6i��'R�+�N#]g?�ˑ��^��g)W>�
�Y�a3�������5����ɰoo���̲�`h� �M�����W�e�K�B,�����p�#L����j�Y��N��Kt�����)����T�?�nk#�-�,6(����W�w9�i���[�n�Ny���/�@���K1,g8��	úќ�q���yi�����m:$F9�#�B��98���bԼ=E�]D��asd�,ӌ��a� ֝��g$x�҇�p��q���?'x.�	`�m���, ���_��/�}P��)nFT �RM���(�)�nEH��.)cƝ<d�
m�:�uy��I6��ɱ�O�آ�NB��e�{���J<ٚm��5�&h�%T-�- ���������$�L�1����^�Ol�N.[��.��و'�9˅��"�?�W�����ц�̓t@7���JB�� �Qכ�pH�|��O��Β-��P*��L[��q3kܓ#��B��OgB�[�/Zp��kE8�mD�`d\�
����S=�����e�p�t`�أr�I3�Ȩ;U�x����ɖϧ�����*�PO���IBE�GV��ze��Ԙoc��F�s���I�-��� �`�o���^[�Q���AI����k����Z���7[�9J���iD}��/�#�]a�#��м��\z������'�1��1�����ϭm���f�/��v"�<��}a���y�b'�.��cԾ�Yȥ���,�����|5� *�j�h�z5R�l���Jk5�͏���U�-�f�N+Wb-��sC(�����H�aU�$[D�g�Y������6���M(Z�� <������V�#��{Zo�����?�|�_���7��+�P�m���jk�V�6�_A�/R6J#�U����J��YD���Yi0���or��yHSik�AK��wXK!�9o"�"�7��>�v��A|��-+��=��a��3��7}hg����W?�	�_h����&�a[k�B�"�$Lx	�u���'=�/�u�|��BO�LFY����ZȈ�V����o��&^�mV�/,S�_,덛�.dNg�Ν�-)�I��۝�e�ML���JW�	ϒވ�	��>No�
��='���l<�b�\�;W��vQ��;��>�6���R�ĝ�g/�bY��1V�-�bKr@=��kum/�K=`V	g�=�s�T��W���d��o^��k�p[	�=��?��vxג{�؎Z�;�/gg��c'輚�
$���@l�Ր��Q��t�R�?+?����٩%�Q��h��0G�T�j�:>�����Gr���7����Vwl�=������;ώ>#�T]��nٜڣ��_��V>hgme���/T<�yJf)S_!�+0ݖ�$P�)�W+��	��n[�&yYCÖb��8�HX9�-��=þT�)&�?�����٣d�N;�ºp�z��B����q���U�,��ا\�p]��J!��)p����I	h(6q�����(w�9���n4�qfA�9��tO������-%���@(�q�b�Q�"���}�Vv�&��P�Ó�u�nj;<9��ވ�� �!��S���z&�������HjYJ�[�N��8��9\(�����nuOs��"���}��{&~A3�����s�ʹ��:6b�m~�Ө���2�,�Q��<͒9~�2�3VK��������Q�f���������ɦU�@ZւpC�����g%m�,��z�7����"'y)��CZbP�.�����[E?t[jnD5�dF��tKK}�8�����\έ�g<���(�iu�=�~� K�^�N~��!eTGX� �A��{�xM�$9�	֡=�@y*O���:�b=�������K����)$f2��<��`$�6+�9����i�h�i��!d��!��I��P���������(�)*�i�]'K�	�t���P����1�g!|��XP
��ے�%�O�h�OH �a� ���7��� �����fO��"X����L�W"������2�7Q#��<�W��$X�T�W24�f�CK,'��@�i@=)~kbe.ݐ1o�GqX������鷘#��G.|#�����n��������/���)oh�V�Pw��b�6���#s�`�FY�.��'�ڨ�	��
�ܴ[��
[u,�4���d&���*�h�O���*�����\����۠���1��3~���]���y_>�z��<.����OF��� ���ǒ�"���Hw�f��#3�����GG��V��p��Ҭ�y��~�OJ�J@�����\�E`pl�a� ��-��q�|6���k���di��Ԝ�Š-F�����9b�є���Ѧ��r�	B�J���e���5�ٖ�4o��i�nx3��؁�Ie�ˏ�\�B�Z�Cn� ��n���?@�h$�STB�-ӱ6���V��H3�?[`��(��cfJ(���F���S����W͚����b3�>B���p@�1�����c�:���~E�Z��E���A=�����1�=�C���w�;;Lx��[J�e�	k2,;�M.����^.���
k(c��^c��tx���T\L"��� ��	�BA6:�\{[13z��M��e�m'3V�[�1��������R�Tl(s�������;�h�����!��0�n!b� �#���ձ�H������f&+�(�l�Ov�����y޳��vQ�mTPdpP�)�_�S��j�mD�W���A�m��1:�S}g�7��č�9�׺Zw�I�:�괐��k�r��/����[`���g����bD��4�A��n�fa��x
�z�(�np9��o��w$�1ъ (O�s���{����X�N�`������"��,�tvk�㛈ͮ����λU%�굩��?�^��B���cI���4�j�YKc�[pK��_�/��N��I��d���2��Q*દ�Y�,�e��O(�;ܦ�HG����:6p�4)�f
$��07+��\p��'�84pH{�6��[�g.M}��L{��3m�
�s\}�Q5e���[s"L�fu�(�o�A4Lt�t~׮g�Q���2u�dO�|Q��Vi�VQޱ�9HN�Wa����K�����@.�<�[�_�G����b�8�p��~��P_s-{��Ĳ�H��Ii�/Zt���|�C�hMs��#�&a��8
�e0�-�T�Iz�� ��a�rH��x��_���#��u��w����ltRr���I=�M�qPiv^T���j�Y�Lڒ�E��Q�������4[Ԍ�A?5?�Y�r��Nwt�ޤ⪶��)�쌒 Y`Gy�7����0�1B�^�w�|"8����Cޮ,t��wKD���9`a9:A8oZJ��+�u�{�ߔ./��l`��,������O9q�6�5 ;�xC�?ߒ2�U_XZ8l�p�IڠMi��;�d��}!bS���O�=jM�ub�ˍč=��}̒�}��oч�UhYj[�j���h��{����{��q��v,����������v���7�r�����]��]��J�!|�@��W$ٶFA��5��.�S^l���Q
�H6@�J������}���G�IW����PqE���"��N�w�;� G���[�׬ g�s젻
�95��*���\��t
Eڙ�qv�_�&��VINSh�*ÅH�=��d�ZC��f���b�`�!��CV�3R�F2D�c�.߹E�C���0��"a�(5�l���+���.^aT�Cw�gU#�h����]���/%7�L�Y�5�g�D���r��嫖d3c+a
4K��޾@���!�G���J����D��~���ȌĜ��䩍��:gX���@��������X1mH*e��8q��2Inp�ī��@?`�P�=m�?n׺R��o`]E��ڮ�H�=AMv� �y(���G/��`�"�lE�h�-��~V��9,��j_�����v�|����39����w_�2?��%�+KP_�)@|�N��V"��j��#ѽ�xL�u���ZglG�wU[t!j������ї�dx^�p�Q�r�%}�y�����*{4���t ���a�[P�{�AT���9D���������`�Z����g[�-��I����\�����s�%�PՁ�E~b������j
��`������0���P��|3�zI�u�R/�f�.��h�-�����n�ճf�?J�Fw���u> h}��L��b�# �~��h���;���h1ԟs
�7�SD�BE������rV�_,�Td� �����[K�L}|��.�� �H�����. ���lf=��k����a��G��t�֞vF�o�L��!��^����+�~�s���s�[b��dH���M����K�7�;�EJ#�yI�yu����":_nY~�Ǭ�g$u�S#����H��G���z��Y��=-�ʖ��U�2�!T���=S���8z���A�q���z0����^����â��ꗧ�S����,��D<�l��[#Z��%k������8�\ɉ�?Y-E*ہ^���P��o�B�")o�l����M�����B��~Edk�alTN����Z�Ù3,��ǖ��Ģ/��^��[6�/>�`._J2z(8x�(u�����R� �J]<7z�@�Ț9�<2(����u��~V�f4������+[W��c�ͶQ�E����k��IO��,cBǲp)�l/�B�0��(*���Z�����[hU�I��1	�K�'V(ɿ�`F�)Ot�t9M<���w�W��  �e!73��ڛÓ^�⛴]�jUP(^�e-��#!V*�a�U�5�ɖi��6-�u8ݸ
u5nxGй���j�q%�x�F\Yz���NwE����T�x[�ëbT7��l)D��Y\��с��4�M�vtgL�o��%��.7(��T�	�O6	t�`O�l?�p|�fc�Ie���R2�tۋ��P+k�� :�����%p.�]�A{N�$x7(�>�kԺ�`ʿ�U����~_l�~4&�
)�v���*�w�64�a4G�w��+{H֙�Z�U��o�w�o��b{U���ϒ���E���8Jf�u}d/�t�� fg'{
�i�k׫�k�����A���T�:L���d��7�*crhǽz+�H̡�l�����}�@+jz���3b���g�B��`�`�^^�a�ZY�Cߵ0L�!u5gi
�J�V[:���E�c<�U8
@���J�j�k	p�2����Ğ�z�je�B��J��l���k"n��cv�h�5ay:�7�s�[sTYf1$��5(�j��M�r3���:qf�W.""F�j
�ys��L�*m�Yr��R�I@J�J�%y@��薟��ĵ}+�`�A^(PSi�&���%���q49.,��x&�tq8Z\p�0X��+�^i��6��q͘��;���E�� m[�Wt@�ʽWj�t��z��KSϼ<�Y��av�u�fQ�a���|�T����3)�E1N�׸������<���Z�۱�qF}Ɯ$f��B�(��N���R��گJ�{ ̩��r!�Yֵ��f��R��A�%��~n�����)Vq���m���X/�j� ��J��WRK�#u�Zku������z�*מJ��LC�.��wp�jpȁ�́1���D:�I0X�X+�@g
��l]h$�����LV��ݷ���������<3���Sm%hY) Z���=�tsI�}�@�C�A������#��I ���?�!�u��Ï"6�ioߞCH>��]��m�q�S M5��h�L���չ�FZ�v�Kvb�H��68��f��҂>-��@NR�cG}�~_�l���_ǋ����[(�-L_w:bnQ����#�2��`�2u �K{M`�o%4�a���lS`ú�H�.��/r��R1��A�3���s9e�*�k�؟`�^�W�|�=�AK{r,1���_8�V3ĳ5Xl7V�
;K�����n6�P�^�U�}$(9��}Q
���N@C��2�Y*G��Stχ����j�(!����je���]�ųc�a8��N <^b|p��a�T6�;c8�s^�wx������g��z�/K4x�>א��w'���L�j{��E��v/�K����X}�)��,����$j.aY�L:�G��xޤ��'d*��ER���G��J+�j��$9�}��y�5�6����8�Y sP��u��'�SS$�ĳ���P`��_9�7���L��T��!J|�*����p]�T�E�Z���3��ܺ��y)�i��W�}Z&��c�Իұ��s�#k�l�e�B�gX����}�([�>�~ϊcxYu����S��x����NO|��zkqe8T��UOf?c3�ĳA�>R�yMm�
i��%Y��YVHa�y�B�h���R#�{�`L�/8!��F��4��;M�/o�Ϙ��� ��~�i��7�w���⽁jy�1®*S۩��m��{V��Ђ��{�U)��?�h�%L������_!I���K�r�坃M��b�����e�\c	zx����"$���aAuiX{Uy%��M��F@DQu3Ɉ��s�v0��;�6������_:v�>6�����a:ש���W+П��|ͷ������t�È
�;p��II����d�R�HH�W*��щ�Z���K��h#o�w���'����&��/�")m'M{�X#�%,�]��v��|�l%�[P�3�Ș�-k��n��}�Ѧi�*WH�ĵhH�G[~����A=���A�4������z�s��,/{R2}�?C�)�o�l�u����V�<��t��ܮ]3���S��I�E��co.�ML�0���q��_��p0����D�o�$)ҋRT��^��0��Nn�-� �Ҁd�4�V%����(mV)a↌�>�d�$0<rdd*���F7��x�}@1��A�;���?AkH��eGٜ����4�57�Y	5�K�)ߣ��<:F�ֽ��kW��>z0M��3!��!`.���~�	�� e��MM=����[�]O�L�3��&������f��qⰨ��7}}��3L螮5��b;8��RxKn��hTbb>󰥎AG�4��,��E��f�ɩ�qV�=#����B�������#y�pĄ¯յ��A�Aq!���E<s�l��L�����z9�O\bI���l��gѦ)��dR|1:�׈ ��A܍�k�8A��%��#ʺ�Wl��⹫F�}�|���~���7�4�q��0�+�}��t���ݔ�{6U���C�#� �hL#�-��nXXdig��L:�9�u@�����#�JƩ��VP��2��sס�6�qY��
K�8ϥ�����~0q��{U��xzw���5m2 ��ZB*�&����FI�;�c���ˆ��z$�B!���X���m��5��	W辠���V����dj�b:ra�gd�D-F�	�ϒ�Mý��&���v��\�FJ8�^
�����Cޮ���T!���$�+�Zj�YvsU��F��������X��n��b�+�����6N�ӵ˨�����ͪ�q���Q�V������g��(�����Ͷ4Gf{�����3ZK�,�l΂��aw�(��pf ��ޢ����(���K��8ڔ�1��]���8Y�iۖU��W�"��v/u�y��M�m��eŒ_yZ�-噷�?CހP����42Y���ΗV�cW�E� r�G�3����낹7��0X��5k3+lP���|���[�l��Ν�QB� ,��#���}�WK����?_y���}�qz62�cLƕ�U�����٠�$h���a\Z$Bf�^�,[���+���Tڕu�1����գ|��sFGF�>>z��W��t��KYU�{I�ÁcpKC��n^�1�혉Ӎ��{����@"z9�2�k����e�U���&�r_�Ĝ�p��k0�j���Y·^ۍS�۳:/�����(E��:0��_���Q�]{ܕXmf�6C�{��_�T�!�������gG4�I<ߴ5S)��M6�$r����d*��r#Q3�E�k/+�5P���Tqf#8�q6:��pO���x�����KB\�
Ih��õ�6�A��9}�ë'I�f@'���:+E�[[r��w�j��V�����Il�_g�Kr�@?�<�#�`�oس�1���x����or��`j=�H����c	n�tK�j���ˑol�PO3������qΊk�%
qʹ �����b|�|�y�#��IѝF�o5؜��3�-�]�4+<������+5��P$��I	+�=����\6��h���=%^�I�pS%�3��0��L)��b?�(+��6Q��n�+� ���;nҏ�d���� ��D�;w�M����/�T2p.{��K�2
��k{���٭��W��jq�YO!���+�j��a�ꎆ܇[�c6���4!���H(g&���X�[��J�p)��LZ*�����ߵdN�K���f�3bZ��"��`���s��8-��N�ߵ;�6�z@#)�
�XD�
iy�:@E��5�.-L�����]���<o��
��Z��PF��TV����:x�S:�W��c	$��B��R��㟛�����8χ��h.vR|!.Ϊ9C�SIã�T���.��ORYΔ]���&i~� |4d͝!�@tyH�z��K�7������<{�C��{H�A{�1�O�s��	y��Q��&ʹ�����C�Ļ�,O��ڂ�8��&6��v�N�ڗ��^<H�X1�L���y�]X1�@�=�qR|��z>�z_�~��E�kb���E� 4�P%�e���h��у[)��H�,3ykO����J�N��6B�$��Y���$�FxL��rL1���`a��xQ�6�er9��R�Ӂ
/�K�k�4�3fd��	`������I���g���b��z;-�^�{�faGۺ�݅ 2;)��~��k���G��^���X�΂��u߽�M{����?d{�5X뢢�����)�����{='OS�g�7��m�+�#�:ZKd�,��\� ��j=��X���\�nwE��H2���!d��K�&�h�ˍS4l�.`�wU�V< �h�i�.wÏӝ��;)d�
�N �e���}]��A��X'�$R �\���<�� f�u5 �2��h�Ǯ���`մ�tJq���q�7�W�"])��8)���ʠI5Jj��OK��0>�C�$peo�A
"r�5�=�Mq�rHb�p[4U`w�BU���}�ǂ3Ef������V���_���j�����TOؤ*��+؉i���v��ں��졾֒�����Y�k��1���gI�|?�h[m�xW�:#OH���է���Q�p�:�a�1���z]��K��f��B ;�~%hM��_����~�={�h�HOJ�T��;�q��6��e�!O�������t2��XD�}Y�{��n�]kj�m�]eU�2
��I�~l߭I>�����|7sޑ$2^���a�6s�U	e�t��Q��9ۢ��#~-����%"��n�
�Z��VpB�%j�;zȠ!Q��M�Ǉ��Peǂ.sNTa*ml
,`#�W����J%���T�����\#�)��[.iơkA O�i�4a��wz
��� �_	è�C�����ɛ�X�{څ�B)����̧x��na޺�KݹG����a�V��*u�16�������9������|wV�&m����b�K$^� �Y6d�z�>=;~���r�z-$a]�P�[�\W���Y��_N��D�i`����A1��L�f.�8r0���	1Q�	��)��~
T��p�s0O7�n�{^�����*�x�'�Hf��<��)�X1�T�s�̗/aˁh)%��^�����%:֞����^���0�7ѭf��>ɒ��lm�@�2�9�<�+U)]1��
��{��|hK�|�3���v5>v[�7g��@<O���c�l�5h��~y$Z�0ռy������B��bg�8풥9�L}�>P �_p�x����*�ϤԿ��盕&w;.f�T`�r�Doi�:��V��9��(Z=$h+B_K��ցj��t	P���8���s��u1?��005��U	�Zޘ.�e�P�9�s)k�͡ !��~���0�=q���%�6�S��eT"�my ` H���4��4s�*�Y�#x�pB�̨�|����'ma}\���H5sw�F��.��@5fgTj=t���DE/_�C���<y�Z<�f�oe�ӛIq��6���h,�w�M�e�!(�n�����d�!�:$0��U�X,�AR�&��"F�CWBv��$f���w��T8�"�����"0�`TM*������l��U
M��Es[���ȂS���w_�j��a�_����-YOʚ ������ m�=�|�L��9L��U�0���B"�ִ|��+��YnP2ΐ�'��E�F�Z�Bs+�&IJ���zk&#!��ɸAb[{B�=��,���j�{�[O/�'϶�ag�GX�7���,,��ܫ^Y��`Z.���`[�'0�  ��\�5�[���ߛ��*L6Tb���Z����9o�A�Q[���^BMU�|w�f<��T�����C^Q� �{��eyGt9�$Nx�E�I�7���Oz3|*� �
�oV�8�%����W�=ax�w1�eE���8ʋK���+��=�} SB�F�jc4r|��S���W;lN]< ���w_~��vbfm�a����+�p��=�$�mS�bG�@&���0o��s�6� ���A��k���Ԯ_S��"�(}�ӫ��`���c�sl��!�%�%��#RHQ.^`>okKM�Q��\n4��xM�U�Ӛ��t͜Yr���մ��o[73��c��qr�S־Qf�:_t!x6�hf3&����9<'�Ҏ~U~!��R�25%�2\@,P!.|%�5�R��ݹWb�̚٢���Jq�C��e.,����rp��[2�3?�I8A溰�Eg5R��#�o��v�]k9Gu$�԰��wޛp&7�H�g�4����9�� ���[�W~͈7�V�B1�fCO$�s�����M/���rq�\l�����R��1�J�����[�c���Jh[�d�#��o\>G'��Ox��~
�?�nu
0I^h�%,�t%�^3��w����=N����̣�f���x�9FaM]G{NGz�lf�O�,:v7/l���w$� ���_ڛ�Oa�k �U�Ǎ��t��
����Ѵsx�n�s\�yհz� l-'
�e!)�ި`� ��iM�{R���jj�!m�&�٘dtb�^�����YyF�HE��X��p��Z��;~(�nh.#�ބH+�\a�r�o>Zx��Yez�E�G�0�qiY��"�y%�\�`Ŭ8<O���ڥ?�.wjO�J��� L?��*4^qbD�-5z�?�ÃO�.%I4wi3{���]�x�q.j���!F��y"z�g�U�cl����i4MB{�s�N�Js14EA`��*n��-����Vq7���������X1��\Zٞ��g�,g�&Y�߲a�ݛc��z����Z�oTqC�>dw'�/�L�ƹ�m�=�K8+s;�L ����h���<��R����a>�X�����A�\ߩ�P�+�����"Ғ��H�E�����N����U�ӛO�M��=��,t�!���*�
���e.i=,Z�P��n�t������x�߲Ɠ���B�>�"�YG��K��������2C��\x�F�&�8^CW~�w#kR5���C|)]����g 4�9�XH.Ӥ�v�~VΑw'ը<�WDD�م��c\,��E �U��D�����bK�'i�p��b��1��i>�'��\��!��^�����+/����gE� ~dWF�m��������F�b�;-���6�铏��K`��模tl�#��$���f�I���qFe'$4���UpǋI��g���Ipן�6 �n��eovBi��T5����B�[ ��p}	�s_���Dz��1�/j�7��ԣ_�R��e1aW�Fd-�b����[�p<$�q�)��}5�0�u�Z�&�?y��=��m�J���hxB�ɠ"��]?�,e6t	w����X��cR �Re��/�T����W��3d[�X|8�)�LJ4Y%rAR�1T���5�R�O�t+�ϓbB��»�g�S���gKU�ͫ�?�*��ZWdi+@��1��A���j���FK��]M��[�4��=E�B��]�iG�	v��VD�\Aoc$	_�ciA�L��q��	�x�M|���/��d*����m���9>���B���O�=��GV�K&(k0�E���<�#�Նd�S�b6�T2����I�+|Hu�d���d�1aHC LnY���]���b9V��a0U.� u�p�8��#w��M���)��G)PG�w�w�W�X7�Bˆ�].�B��ԍ0���0��P�)��i�b��0�[�D6���b�έ.���]�7�@l��X�Z���h�~�r��y)�h�����8�A�Z>;z;�v��� u/7`����V:���P�U�t9�;m(�q�~�t�ijX��;�Y�)'f��
��\L]�\h�X��z����u��ha�o
�����9��?D�p6Sk]|��J|ĻO5��7n{�mY���<���i��&���	P�׊�R�j"��ʀ�gU?"=�?�Oz�����ĥw�����C��7�@Eۙ8��.�s<�i3���l��"$_c�8��ŅA_�I���[�T�� �T��{�1I��(�U��:�tX���1#z�Զo��Q�1L�����WEx[}c<�&S�1�ׂ�V� �d���P������0�hO�dO7��ڭ��Zfp�2�l`��OB5�$��\z�$WLwJ�������&m���Ĝ�]᱒�P�,�*{�w�R�C��'s�ԡ����E��T����*6ak�E���E��% ����K(go���s2����Op�^�r>���Bx:H���*aR�Y���s�\�BBFO��L����'���P=��b�ĳ��/��pQ�Z��vC((��r��	�������R9�f�����|�絏�H��g�`��Mp��w+������m��s�~<��[�-,�ogj��	q~�O48�y�/�R�|�?HF�7ә�3��3*sx�-��&n�_��^�lY�E�~1_K�.���e@C�FrsY\��hE��N޲��V��xp�3��CJ���������[Ħl��� �b���&���2��Ԝ�(��CX�ܩ�ZD���`rdN�qAb��=<�2%���օY)����Y�u�ێZ�_DHx�v<��=�;d�7B���˥ùd��h��T����b$ ��N3SĜ56�
���%8a@�<���2�����R�m�����a)��
��çN����jҙi���j7d�Rl���D�޲�����P�^�>��bԣ��3�?>M���VT)�MUI9�)W��P��(�^��c����,Q��:�%<f�Tl��J���Т��9tZ����H�-~|Ș)/H�y�j��]Λ"R񨔭vU��Μk����r�"IZ��n��ߧT�Շ�����gU�Λ,ML;ܦ�|����)W�>�!uQ�]pip��J�W�q�M��3Tǆn�����.�=�DIM�}��ܟ\̩3�/^���	�+�q}��q����Eo�ͽ�C���T���V�2�ˏ�n���]�[4�M�F]�F�BK}�]z�*����O��Ȗr�^�O�w)��o`���̡dx����_,9K���Y,�?�᧔.BH����Qq�����|`�"_��(I�����K�&�&��~L���Bưp5�fC��/� �-f�s	;O�������N�I϶�����6��,#�=W�`3и x��x4�V�:�r�mw�Y��L�ߢ/|��i1��ɿ(�c�}�Ä��w}8�����Q�/��/���6�Y\��Z(�V1�����ls8����"�b�+�˻���J�4����br���$�qj�w�&�~C&WpU�Mm�L�lO���&J������eD�z�#ué�0�����<qJ;"]�X)�MqՂkfҝ�ƈ���1Ք����	�]<B�;��TFpx^DM@x��8��م�r9w���K����[�rA�]c�Ɉ�Xu7hS�A�r��I�A$��&��)p_��`@�' ���5`��R�S��q�G���Y�d�g�4��~c@�VZ�����Q�x���$�|�Մc �����	��' j����2���f^-r[&P5}�Ƥ`�Y@_�;����t-q��{,kL|�y�?�4�/jJ�j'p8��7BPQ ���٪v ĄI_<
M޼����]�jh�M��-Kw:= 1�	��b�L|����nl0ݚ�0��:�-�C��nU�8^�u���ծF��߹���`w�a�T��Ѹ��m5h��Y �s�8��K��͞k�Y�6���;+:�����W�5��g^��^�HA'����!��z�}�P�;�B��k��6�)���$;��-�3a���7��w�ݧ��y�M�O�Ũ8��]<kD�xΨ��;��y$Ǯj�*��fF�n/	��noz�+�3}y�)J2����MN��J��W�BJ\��=���%`�yc{��iRפ���C������AhUT��KP�Ƚ%�؝�H�Nm���r����&X�{��������������W�4�%8��=��+�x�4^����e�*���<X�����;��,�8�
�L�������3޶�q�>�?q�6J?���W3�Rn�vD���5� R_H�t�;�	b&� ���i��l.��M�ڦ��J^��eme�~�v�A�&^AbH��}�/_���5�"�2՜�i5�a�HQJgB�8<*bxY?e�q�B�V�[kz�~�?�� �m���?����X5�/Ξ��:У�M�n9flv�MM���ւ�З�r��t�c�m�0^��D�����1(��|2�4�t}�$a֙ѿ���
�d/ϥ�&B�)uo��*W[SE�m�)N�H���H��:�O_)�[���w�ז���bh�C!�.�=3����(��s���SFy�s�����d����{Q�L�N������[3�ٰG��<�s�)��>(��Y�RM���˦T�G4E�G��-�!�>f�E��C���*h=1&ǃ����n���E��\�*�i"�;����d���0�b�#�T��tI��;E���B��%�����,���y��Ƭ{3�ŵ+Wk��� ���г1��i�C�T�&5�է)t �@-d_䦕B�ֺ>����"��|�Ϭ�����p��	��0��p��"�|��m1*ϗ�	j�;��<������J�{R�ICM�ᣈϽ��'ŋ��.�5��S��*E�,��<+���т�:�GQsW
9p�cY�p�:��/�ٟU���ڸpcKN�gK����r��]|�|A�x�@xjB�!��_��n�ޖe�����yұ��B�K�X�V5x��V�Z�$hreP�7�J��p�I[H�����&~T08�����OHV��),�$��bzp �a����栥��ɲ�g/���w�x ��g����9���^���^W|�8�-!��3J�x*����fʳ�t#+H�zEدRI��m��];_�6ߐi5�����y޸�Ը]�7�ƺwR�@��r��L���5p��fe��f�X�f��A!�vQ	@�z�c�@Q�}����3:Z�0�r(���/��sq`�1��)�;�`���/�?!]���7��(a8\֔����LD�����|ꭺ�h\��=��E�p��q7����4�a��,Թim B����A�e��&<���^#�:U+o<־:׼7~BEy����"�ϵ�*L��#ʜ��^��R8J�$$o&љ}��j�Z��CF/\(V}�)�����w?����+f�Q��{���C�QN՟tO.��p�q\zg���c��Lǧ��Z{<�kz��厲?˥*�&~�7RS�G�8��bVF�j���H�l���'*�����z�hbiO�<�6�5xG�K��xrX.�YPx�/7�yY�����
�(���Bv?�6�(��l�aψe��u?�2&�mu�M�������4i��}֘u�
��8�y�[���&���g�b -����T4IUP�d*��6���D�t��V후uSY�7e~��<1�p�c��L�*�����7DS��W��2T�����U��mCx��̨���?By�~\M�q��5���|����ת�M&T�eʳ�^����zj�	�g��I�ρ�r&Ho�@4]v�楐ÂGD�����A$�K�ϯ�:>l�5F_�/�^|{v�$��Y���>><�}#�Y���U�r~�ww�g@��=m�����^%]� g�zOl��	�LfPE�s�b����0�<y}��{h+~�s8Nܪ՗1�v���*s�rP�e��j�tn�]�$�9�b�Y��k��m�	�'�m`,l�j��i�F�e���U�C�ia���K)7��+\z��yQ��>W���J�Y���{�9dT���W��<��H5�IV����e>�cu�S�/h��&u��Ѳ����'c�|-W���@�V�R3��![j���i���Y˙�U�Z��ә2D� ��	����KL��l�$c�$����g�b9^�2��C�����ו�	���j8t�ĸ箟�w��F�'��ϊ��>f�v���b�kg��7YV�$@		1���X��t���i�~��(]1w5���Gp��`�+U��ַ��I�k�f�N�~Vj��v�A�~'I	1����2���td���u�>i��e�����jH�SQ4;�:��J�~�/��Kϗ��@Z�؃g�o��AD��Eۀ�q?��a���[1���Ֆ~U���z���:,;ď#ɏ;��a�a�^N��}�g�<�r��[�/+�uY}�.�Y����w[ ��8fS7G�|�м�)����X�`��)�L�7��ؼ����WF��V 	)7�`�r�B�;�a�n��!��)�\뵞���;����|c� �NW����ڑV���&UD�G�� E�JD�7�}�{ڞ�(��r��bcy��;��ѐ�&�oM (XS\���@�B�*|��_�9�X�5ŧ䦌g~^	�w�쨺6dq�<6�Gε!8�#UD۱�v�4��%��/aa^�ZS�B%��t��ڄ��1�*�P��)Xl=�e?�owl�%����O0ve��
�삗Q\��O$l��m����;�Bo)����h_�C>���*FZ2 ɕi�Kh��D~Xկ]����YIFk�޸�Q<%6��òψ��r��>d脗'm��� e$�Y�♬�t��^ ���_�F��?x�>��C�f���؜�yD`�Pc�Y�h����4����p���s�rȫ�D��(�qԘ�`�5i&������#�^��10~&���6��A�e�ϊ2��.����[��\O#�X8��n-���H90�{�ať�|v��6cޡ��PA����eE�=��R�D|�5�ly��"��� �{/�v��TV'��+1�_#���#��m�3מ	׼��hj<mC��l����4��8�Α���;ف�=�*���-��G�e_���;�� ��gd��>��`��5=9�J�z
��.ߡ�h9��m���͘?1� �~���@j&����p[��  ;�M5v/,t�R�-L62��}�jq���P�랖�u���8e.{g��\�7Y��mt? )rk�4I��Kg���.��ۤ�Be�C%�k�Gz48�8@Hza���������d{���֐��D��	}�Ǧ�d��5���t훒�ܤ �������~�h����Xl�mK��ʃ��^��z[��I �Nv?c�Ԫ�j�
�z~"�7�%vΆ�O�G ����i�4&���P^gP����]���a���j|����i����̰��k�
s!�#��SRq����"S�9�*�F�mO3�+��Ԣ6��W���n�Գn�ꄡhʣ�wԒ����=��<�6��ͳ[I��NvT���m���~&??+Ҹ�����Z�/��m �:��T����#r%����X1����V���'���kg��/C�%��|F��I�3�2�I�Y�?Y���"�����2p�qC�t���-Y���d4���6�~�^{����^A(�F�#<6���������ua^Rk�?m��F��_�*Q�z�<�#�ţ������m.}J��9�_,4��7�p(��z��s<0�/�b�*����# ���`�'%~6�6w/�*�|�aG�m��_GT'��MT��<�gJ�K��e���9���*i/�T>��$=��E=U�9O��ཏf^��}7��1�E�W(A�8����bs�UC�V��N��D��g4w�����UW	m��,��nM,g��Z��3�X��ͷ�7Y����*�)�I�
|��~��L,�9�^���7+^�h]�{ �l�@9���J\;(����Qb���#9���yS�>\X;&w���O:o:a�ƒKe+�	����Q!���{'�N=OX����5d,����W|���w,��igqI|���q��.�����%I��,w�1�A���GDAe��{g��x���r�V��HΗS��tfD�Ŕ`�}9�̕�3	�΄r���$��`�I��D�7/��$��}�H�T�fSDSc�Ӳ����#�9�z��߯#g���g*3t��.
��F/l�,��C��K��|�w�ԓ�f�C��ӵ����T�'� >�R�c��m�2em�4#��s>���2�v��!D7{ ��#��U��\ɝf�'u�y+���hwlD$?�xM�u+�'D�og|�ޫ3�ƺ�!,ۖmrAZK\���9�^�"-�ܧW�'�T����v�@h�"��~me�L���{J��6����$�?P8)��}���ό�4�zᡩ�n��x���LL�_j�`O�|o\k���X���>�%��ܿ���Z/��F��32��i%�"�m�e���}LW���i{�H�`p*���<�>&=�A�|�(�g��P_���^ʊxA� ^e<8�l/����Tj��<weZ��O1��bZ¦�&�z�R�C/q�2BP�D~�ǿ��<$�`�F�zsU�.l(�ZXB`�'���՜ @ʅ3�,S�m?�������W�6
=^֞��s��a[�Ta��a%�"-#����'�zǕ�E��T�!a3�[�̽A�N1"&�r��
&:�2���0G��ں��Bꄢ�Z�Vbr	o+Y�����a����9C�lO%����4�8�@��A��Q2��;��L�ݮ��!$�&�CΜ�i���H�"����-l���h���BC�Kv�f�	��q��0��+��B"l
�`�QJ���T��m1f
�b/����ި�,������nP�:���X*5�P��k(�&�I\ݹ�\?,
�N�B��ri�GK�:Ŀ�����[��z���A�.1c�@�H�#��n����\�ݬ���������hSߵv�|n���;Y_LFOi�)��e�k����/#��Ӿ����2����*�=�o��E�=l�x4�����9"/�i�HG���؎�a��8�P��=%�����gy���}�AR$tR�;�N��>��W����-/����^���2���A��&��E�_A���{-:(��B䨒����'{q~�M�f~������yc�h�A<c~/����X[�f�Pժ��L?�Aw�7Px��G���Uj�������g`Y�����"[	 F>�����\�*y��B���j�2��+H{��ʒ5�Ou��I�뢐�9�)�w)����Qg�B֟�=q��B�J5D�f'<����ɿJy�_��գ���?>����<���wLh2��9~��y��*��{�G��f�p����M�\���\�޳-��O���,8�f�ʋ����7���.����q����ObC�s(����aE	y�~�{�p�q��b	�$2�5�h����Î���Nі@����!+���h���m���J܉'� ߇*��:�g���?�BĐ�|�����Ĩ?���XeH��:Rx�`��s$U��4a�C�
�=�H�yy���t�k��>?�ǯG-bG���zuzQ.�5�����U�ָ���A2c��ϫg�ތ��}�3�L����y~1[9裮m�-�nKr��;�K�����dz3_�=8���J��=���Jq��$��"MJ8��qI"h��옣�H�!���Xi*~j<|��E�w��E
�D�_W���y�bf��*`V�@6�qz��c�a��Plvc� �	K�C��ç�X1uH)��R�8�î�v�'0a9GJ���4��:��㖓\c�>_��C�ߘ��/^DbҔ�t���s��Ab��ot���=JsК:���1�c�Jdd<H���)w
����P�&���n�|?��`�C�YI�uD¥�h�
~�Qِ�iȰŞ�h����d����q�N�5��'*&U�S;8�ggŠG���(�:�:;|ṳB�o�s����0YK�?Mw�]�e�\=��Ok9Hͳ���nr�����-Ƌ�o�g�#��秒$+�U6{H�Z�m\#J��4m�z\��U��.k}l���ߎԛ����ɿ	����jan���t���}��t�&�o/�ҽM5��XSߔi�����-Ûo�ΝA�q���O��D�'�MQ!�}[���ƩsY�x��Xd\hI'��f��wg�*x�4z�%��x������8R�B)T΃�w|Yɶ��h��0����K� Y���|�#+	�v^�?ޕ��xW9�{�
+ӿ�d�iSA�>��O����G��LF�'Bk��b辰����޼�~gNʎ�1�?Q���G�����҄�)�LV��?��SA))~����/�2�G�,�����Dq(2ɯ �� G²J�K�:}� ���O¾�>�Շ����K�ʡ�}ka��7�@������ w�
l�IۑV�м��.��>��� ���L"�BSs�'D|�B/�s�`���x��!�q&�q��5=�[>�5�7c�-�k�E�E8J덋.k��]�ЈǛ.����<0..XӲ	���8ã��A��5��G�!l0���,�0����z>�{a�T�~o���V�/c�q���n��g���N��4s
.Q;�T�*��[jq�ͥ8��<�������r%�sW>9�`_o�`)�:[�J�/���H���&i�&��*�H��$+j]��1Q���-���$��:�nu4��m2���[s������#Lϻ�)���W�\J���;�\�5�H�v�ּ3�[[A4W�"��*�7��x�(iyj�rh�sPa�=M���~�E7�](�x�*0����a{�4���"�R�2��pn�GԱ\�����3B!��HGLs�Q��=���fd��g��1!]��C|��:�²�����ڦm9<$�l�ΪY�{{�
��K�0�-�'�ţ�cn2ŋ%ea����
��[�KeI�����Pļ�tet�D t/Ҏg����#�a��F��`L(�d�"%@J�E\`s���̏>�|��i����\��+�����m�}3
`��Ch6D��Ul�G4�T��j3V-=���'���a��|*�6D��1Qt��]$��P�A�s%O�s�p�%�~C
!ɩ9�N�؄3
B��z�V��w[T/儺��v�fWHT�7��~�_F����U=}��]\�[��������^đw	z�/����́�W+��9G�{L�����h̢^a�e�LA4VHh%,���X��[������4f_��X�|�����U�b��62\z�SF��5�%#Ao4�@�^8�>F�=�X���A���ß[�n�g*W̥�@M_Ѳ��sxW ����cf��Z{��}���Mw�Yp{NtmmD�B�]9���np�p��q�_:�If��1��>�.�D]�tl��:��'@8]�1�;ia���\�y�+�D�E֐Z]�*��UzLX�x��L�sv#�/�|�C�8,��s�Ɇ�|�1����+��V�༫7��8[
�A�6c�=�I��CB�p�WC�H�M����)pv����q.9i��H�r4�8k�C6$��T�lB��sU�ӽP����y-N0�%�ʹxy��2���#B:yD�p�{4O�h��U�Jgy�aJ����!�a`�ho�a��P*�;E'�z���������&5��K]ҥY%���uZuM�����yN`=�
]j%'�|	/���0h���G�a�PR��X����څ|7S�؎e��MM����'א�;�#��$�ݳX�g�V�� X/Y�Q��C2a*��qt�X}���ƌk-M�W�(梡���3hl6�7����N��x��|u�abK���f���~U��H�A�� *$:|7��#�5[���&���$��;7'���Ġ	�::�=�ZK�����~}
g(?���+h���{��=+��ۿ`�Y�͝h�u���ZY\4ʭ�V*��L��U�~����aJ�A��a6%���wK�d�qn�[���*�Sp�o��R4icȡ�=COP�Bk`mO�<����^9�71h�Ll�O�:��K���X:l������C�|�񓙘=��X�w)�!N{D���$8ֳc� ��:�Xf�L�)<�i?q�P& ���~�u�e{�+��t��m59;]%k�&Lk��Pi���_i���\Ϡ����[�����P�8Y���GGW�U�|Q������HO���7=��{��.o�����
��Z�2ܚ�j����`���O�m�h��v�(s��,v�%�@�~�*�	���"|Ìt��L���g�b���z����tl��0��u��@���*uCu%�gH+i?�=��!��C�e��q�ɏ|N*����i��a0�o_93Hzj�G�����Y�T@͜,���ec߻ $�)h�KGf��s(퓦�M�L�E���+V�I9D;%���z�(�P�G�J�Y����Ӫ�yES����ͿُA���m�C��\���z.Pc�����w�1w��Tl{IOW���X��k�Eܣ5�|�e+��"�&�H�Tn�!s�}�Y]%Ōg(vb�0��'�tu8ۄmn��h|~Ǧ}/��������K�Ҧf��(]gy�f�>�?a����`a'7a����/���U���#O�%��iWBX��n~�CoP� ��(�g��[ڽ�1��b��Ĳ�}:\�RUI1�Y��]���n{�n:"d���W/8��x⼳}6H��,v!��5s�o�_��fw�=4Ub:�Z���E���8�����	$$C	�DƦ�sr\V�/�i��=�US�(�<�*�\�����zs�O��^��_��9V�� �J�����
�~�(�S4�g���34�$����͹���t;Yv�>�EG����@=�u�(`R�����$�rnG��~������=���3%��0�j���z-e: MD��t2�����D�Ӕ-)~��l���,�q�#��=k���3>`p�o��>�>@�Pu/��0�P�8�8���c����V�k}=�Mx2¾[�����(�0�ׅ%�1�G�u�D`K5���Ȫ�k��޹%��Iǻ��8��Lb��I��䥅帖~XX�hv�YJ�%B4%'n?�~��,r�a��T������� 	3�6�ƥ���	}��V͛��hX����l&�{ @#msp�^l�E/�~*�`�@�$`��euH��GUie߭� bk6d�����'b7�{�Jm�F\	Ж�g�;�*k���Q\�e�ޕ�z�S��c�QFmz\�l�XI0[���xi���-�C�8Y�e��JA\�]w77����*2^�߶6�,H*��ނ٤�*i{6+|�%�[�kŲ��8�%l�����*���C�9�[F-n��˔5U�qvcq�$4��!϶�y��th4���\%/Q�y~��r��Q,��E�|k|x�s�Z�uF�l�Sg��mg�P�K���pXK�j�
��6�0/Y��Y��z�L׭�%)31t�Yh���q�^�ڗ�$���J����p>�W���Q��t�Q4�������y�h:C�N�<4�B��9>�����Z�x��188c
s>h�'\���"���r�e�r�D���N��q�0?s�a=�Q�x\���M�!�4�i���zW{�Ye;X��6�@�-��%,3(�J޿�n���KU���2���tƮ�^Fz=���G
7�W��r�~�kf5r$�E5|�	�WTUi�9�ҧP�]�<I[�2�h�D<~E��\UB�@�k8mӥ��,R�ǲ@~��$�S�WZ�ݓ�?fW������;��"�Q��W����g��A.�ڣ6ۿp��7����k(�M��FS�˙jQ$�����RTѮ��޴3'��C���8�L�n������Бe�%5�P&\3��m�|�V��2���dl��jy��,�٥}R����d$P�ϕ-��+4ה3�QE����>
�a�8��=��Տ2��rm��t4�3�T�3����a�Eu]oJn�)F
ۇ����{��_�.�?���S����A
M�4N�x=[������~�4���V���k7�2tt����9�9.ٗ�G�^c?�6hW�C{
g:�����"�:~���i=#�NPNq�;���?ƪb5�돋�ll���ge��;��u�iζ'nWg�.9�$K��r����{z*b.5Q�%t�`�9`=�0���%>]�)�ߛX�EM��gȆ�񄡩'�Y�o�^��^���cie]'��sz<�e/Co�BޘK%C^r�kz!�>���j�A�DeD��9�ޟ߻f��C���Ⲉ����H&�H)�c;�|	�J�����&I䁢�����5�o���
�Zn���(������S�I���L91�	#ks�]Ň����2+.ң�q��; T�����~��I�a	�%�&9���`�h�+����N�E�m�и.��s��B��\�\�T�>:Mz6� [���9��V��0b��y_1t�̐�H�vk��d>^�L��2��>Nm���4.ϾA.l~���L6T�QF�g#����kĳ6Y����+ݶ�ԥ(P(�2&�\�u���6-c�xgɷ�>���I\�0���:�}������W3�{|+Gbe�� 5)O;Kf�h�k�Qa��|pQa���`I<�	ģQ�M%T;�g��fO�8�]�F���?;�}���V{��IS�<G�ho�ۜ�8~c���D��;O�9(���(��W66�p��. ��1V���e�X�hH�%f~�͔��[dE�2�%��9�;Y���fp��V(h���O¨-�4	�տ��B/�
i��r����y9-�];�3�09q�lv	�9�����.�C�����; 3���>���>�,>��s*�u�S��ZM.�������c&�5��h���%�9�Y"EU�}~6��(���{ �^�z�]��86�"�9��P:֛�J�lDrx�j[����!��둢@#���o�g>�EQ6�K1�
�c瞟�
P�Uצ�t��>+��c��eSzp���w/����^8������G[��^"Q|:뜑\��2�<�9jMzB8�,����~O�̡�s`H�
o��k1�@-����a?r�}��-�aZ�A��Y�L2#�`TY�{{>0����ؗU#V����CU�ň�H�x$�S>��j�^,��T��G��0{zR�h*<o�VQ����q�0x+�HR7�Z�O1��;�y���ُ�����'9�2�ߍ,e�*��? ݮy�o}�
!߆:gOMf+0/�����XJ.^�űx����~l���7��܂ʌ-S�M���/�EU�	��esks:0�.ym�OR5�m�Y�aɁ����O"��a��3q��U��䱃�r�c�
F��a�Ȥ#�w�t�*Ӑ%�(�V�g��m���J�A'C���6��͌eV�!�O�`Zs�{N}z�̾�P�?���))���?��4�C�Jv��)�?Y�}(UK��^ij�˞�s�ȒJ�̵q����8��h���L�����~�+�v���Y��,���|�|޽ܤ]a�+f�� �"���/�h�i�$#$��N���p�,\���X��(�%]���ϴs�_C8�/��	�ȓiw~���!lL������������a�1yb@xoE~k�0�첸Kg�� �m	��v*��0��m�w�N�|�p�S� ��61zD
�K��
���㍆F���a�w������;nzx�y� @�-l[˄�u�L(�&L�A�s~ͥ�e�E�(�;w�v���/"�	e����-��3�][���i�_�O|�}�ӛ� �&ɂi,���~U�jZ��j�
���%J�]��߻#N@WP$Ǒ�gӰ��*& ��E\�O���Ͽ���U���I�O�BN/p�j)�Ur�lN����$�K�t�>�FG��vt��W�3 g���Ҽ��L��fk��9��6�P0��1�^Kro��F��'�w��U�|�k� �����6-;&�^��U�0����X��ʚ
Ȅ!{y�᎟��n��<�sh�%2��p �E�
�Qr�]耫!�l'l,ha����y�:��Q�*�ޞU�Z}�o�S4sJ����yƚ�o�H�@y2��"��tB�-�v�wZ2׍�F;��-^q(�v�4��xe�=i��\��4����$��	����G�RaA�*M��zQ�2�	9܆�V�>�H#�N���������� ����8F)Y���[�?�#;S��-X��r�z��]�]�p�ݛ"�]��H��vYۉ�"_hU�~n���1��R�r���W�5��j~;� S�e���QV�3G�t�s��CY� ;��P��=�z����[;�5��7�}�4'FE%���遡����'���i����@�-�h=0֤_3�[�`���iW�����j/�B��ّ�OYnP�>Zn����X�bj�`���R�o�b��vynU�{R����<NlNy�w�7\exi����9h�:�j`;�����xy���W	��	W�eU���<� �͚�!�p�6L�	���kty"*�)T�t�i���{���XS���p=A	��[.��8�O�H��^����`,Z;�U��n��e���kx�m7� �Ō���Ku>����̽O���"��%��=�A��H��(òu����E�3�v��D2		�2��%���K�>�L?
��FB�o��v.���f�f#'m�թ������zp�s�ŕ��e��h�	��v���`cQ�%N�M���N���7CђlW��T�z�:��j�	�ǖ�M����I_��^#�g�N�8�C
z�o<����b��!��V,�@6�4��P����7@S�����0�����.sU��x��t�K��L8m�P^a3�'2���գk�zxR|f.�����@��y��=>̯�Zv�[zd�����Ê�dY�ɾG+ev�e��-8,G�Pǰ]�X|�ba����[7jVd!S}�z�_A�Ň�Cs�Fe���{IN��Ȃӫ�碑M����O�V��9�MX'$J�y �ɐ�e�l�v�}ϨX������C��L��E)+9sñ5��S�lXl~�A�Mƽ��F�O��4�d��@�h8|gqzW��W���ҽ��J�	�A���� $H�����p�P�&�7t�a�%z�L���&�r�k]t(Pc1�\���v(��]�ϱa�+�H�zP^��mY�fM�J��筀�Z�w7�`��LB�J������y37T�2��]��L$��զ4��gt��}�=m�}�Q�|С(���u�$s5O2�WJ��N���pͭ�/�+�n���&i�J���Y����N��eyL_�K�%����e�$U���h��A�M~{C쭾/}���0�X9[/I�U$��P��d�6�;��O�L6�3k��C�LӸ$�s[����Թ�^K�W:�`�5KO�8����� �x�Ϸ��pȰ���H[�:�Ċ�9`5���T�!gH!Z�4�3�&w�5dJ��B� k�T�z �8�2_�QU�r��r�3Y����m��S)^����u��M��;Do�%�~:�:K�"�EcV�:����Q��n���#�����e����V��IO��jG9���F� a���5��N1�w�g���D�3�6�p$���X.��jH�k��=��!�7.M���?LP^�xc��,���jv`ѫb!�(4	z��m�O[�ܕ���y��ؔ��f��-�C�_��z;c�a�]��Va�2m����;^+�Y�h�%�#Y/�ӳ��SDߐ���.d��ǸiJv�%kj0��S�H$@*FZ�~=n�W <$��;�:���F]0E�2�p����wƫ��7z��d�2U~�]3���P����u�_��XU=�l�_�f��Ϲu�R��{��)�2^�ۗ@M9�T꒕=	h�I�2�^��c��p�N�mO�.�XF]C���s��L�b�L�/==�h�f��pO˨��С�j|E�O|WG��M���=�a�r�4�"��$t,�׿�X�O8��~�M*�<��K�3�DM|b"ń��6�q߫��*��5(.���c62�!<e!��<�iyT?�v�����2�l�{m�_�O�@�b��`�Ù<~�1�Q��/�ZM��:��W-]SC��o@۲9�.�������>i�(��ۈ,��� ����5������s|JNa��.đ�eI侚��~d5az�a���d���Me�t.�;;��e5�F�����G�4V�#F?a��X�+�AIDh����
���=���.������UM�c���j���‒�<_�ˢ���M)�*��� ��p���{�~fȂ&�VA�h:��E�3>[����
�#��E�m�V��ۗ�.���ot�>ݰ���(NB
j}��`1do����_� �4��v�^�3q��PbAr�qWf@�M���`]���Rz/u �%�T6-]�X
D\�^O�#?�,֘quY�"��B��ґv��{�儡v/)_����r�����E$�$�@��"�|N�ƚ�2 ]g�90��6���衍�+�H�|�0���Ϸӷ7HF���I�����U��a��Y��X�gP���h��)FI��(�WD ��9]@FR`���c�z+�{�{88��H�BA��x ̉��5 ��E��tL1]���'����l˱��[�h��=�Z,|L�hdI�Je�X�=��t1M9�Hh��ٰ�8��2��T��3Ow��'W�� �	>N-��mrn�.AW�!�50"��Q��uјkҢ��=�%�j��C[R���@�	&�#ݔd��;��#fO�s�\�T��4��T�r5!+�jxd�ʮ4 �
v�ל���������7sР̳���{��D�hA/l�$?�+%7�(�	=� �th_�Y^����C�I�Ou������ h���`�串�/5~�nx%a��o�RrP.��ݺ�e�ba�$E,���F�n{Fdy�y8����z6���Mt���:lTiMz�j2ض�'����Y,��*.Z����.�G���M���S�Y���W����n+��bBD�a	�}�@r��$<I7ْHS�����pb�.�b�� \�z���u�2�퉔F��x�e�D�/|�ΰ�X����^wY?	�r�b& [�)dӫ]��X���T6��8uߕSwI�V0��լ����~��=F�u#�n�&�B���̧S�e-���
c�O�xj�C�����wRA3�����B�D�kd��]�'�!H���o?��r����5���z
�W��D�)%���L;�����}]�`|�z_��%S��p,��#�E	=��F�XBqS�bX�d2���G�/�*����6�ϙz�.]���CN��p, �8�"F�ǣ�/3��h��·��|�Wγʅ� ��/+[��7�0�k��$�Q�"i5�0�pQeS6��"LA�w��l�v�!e���-*��#���-�����/?T<Y8��CO(�q����-�/�-6��"�v|G��`%h5$_���7��{]%�<DT)S��w35w�hC�"8�9�m�P.��I��Q�O$�b�x4R��YƑ���b�4��Rډ�]�Ujh�6?
�zy���U��#��6&�V�n�r�s���g������%���T�b+��Ʃ!W��,S�g�1USu���܎x:�Y��~1ó8�3�ֶ��Y�2���eno��1�.�(3������#�EC"���;ٍ���C���cV�w4�}� 1�qC��A8�1:I�k����^[8��`>�`ʗ8=|�|�J�I-\���)�RR\7[�RHt��L��Vʏ�ڍ!|���}�CR��h����%/�6D{Ϣ�Cv�<f�87A�@n�e���*ݿQg��ˠT+A(�h5�$礑��J�у��M�?���Z}�D�]��q���9���A8(�u��k���b�����P�H����$*�s�%ݛ� �fA6z�t6�\������ymof=	� d��I���h�IA%#�X�?9P�)g��%1f�ު&	�^��u��B�Wri��lDW��k�2���V.@�� _�.
�� ��ɡE��rxa\
�޶��2��qE�K
�g咡q����z��\��~W���x�r�0�r��Y�wpEct�MI��Gڱ֘Yov���`Y����.]����9�8M&E��U����X~ڍ�x�t� 	�WI5�Kl�.����^��N��'J)���\�GH����Dm{�?<�t:��)����#��Q�^�w�����lg�R9�\��	�0w���`�Z��;9Հ.�W�7����
#�@˕��Ӑ��&=}��Z�t<\�s�~�\ �^z0�Ic8A�"g�#�vfSB�� �����(�έ�ڤ&��#�� �����A��5s]+�P��Bmm�2#l��^�R���`���3���2�)��0�n�LQ.hG;(O�&��u8y�'J/yE�����0=N�;nu�̿�<{%Ϣ�fӝ��Q�5o�އ��{L2�����^�US��Y)��;�Q9+�����GS�|�9�a���r���9�Z��S��*�6m-"�\p�#|4Kq
c��ւ���);����[���%� RWkw��	��=�s6C�P�˰��_ڊ�7ZQv�N@�d�.�������W׹.9V��!�ϾBU��0\Ey3�0�"���"(����F�D9��ZNԵ\$�R�aX_^���Ά�'�0>�p�͛��@Q�q��e�0�=���P� ��R�"+o�W�m��CP�IgD+#�M��.0������K��UB���3S!�0�Lj����9���Ĥ��B:`��v��ʢ�����p�@Bs;�c�v��vuq���d��}�#�SɆ���E|&Ĩ�,.Bv�E|y,��5J�yD���p�Z��c3{w�]��[~ �V.1�`Vw8������?�6���z7�/_���c�s��յ�'���G�)W �����������w>iJ��R:'�"�Z=d�ظ�>�@#��&S��A�&��c�?����^�:�	K���<�w܁ܭv��n���,
���ߊ-������.�"�X_"�0SUrc�	7J��1�����5g����Y��G�ƈ8�M�UnB���м�����A�%,��m:�.�՜�Sf���W�b�t��Qg��@�����������S	 ��ƣ,f�m =���/�Y��/J�һ���	|`�3Z�VDͅ7S� �ˤ����V��2���u�[�vV�yFS���R��)"���WxE�1c��7ǐ�X߂^E�v;h�����.ڵ��]���I�����^�?��I�j�� �Y�|�d���m��C��z\"�Q?�C�R�Ơ�E'v�E~�%�8m-;��wat�jQ�Byq�'V��8��}�I��sW��q�%5SV�zӾ�Dxr���@�~��0H� �h){�)=�j�aB%yK����g��$�_+�ʄ0�Zc���?Lb��7�O�Urh��spY��B�W,L������t~�x�K���M�N8���@e�oN�U�7[-�-Ш�N]� ��#��3��R1�\[|�=���3�s����'��g)�x���#ڸ�]��'"m�b��u@Oȡ{\�P��Q�����v)mLfs�*�� *��7g�jnU|�o��{�Wd����3+��n�/>=>� �k B�I*�����4њ٤1rZMu<�ܛ�6�ƹ���[��$�_NZ��u���]��q�����He��c|z[�|��I��^}��O��DM#ڟ�z�]-N�Y�:���J�yo�5�I�: ��<�e�n��:N 8��8���c�V
0�Y�ͥj�ueK��c�z�	.��Aat��!�/	L*~��!������:��	�j�O�5s��FuZ�P=���z�2������3�R/�Z+��rH��ՅM��>p��H
<�?Yh,�db�U�"��@�VW6����c����0N��JE��J���jz��ԹĆ�"�>q�� ����td���a^�l���d�*8�����P{�Σ��a�!N
���8�É-�N�CX!Ĝ�*�[Y��7�
����` ��#�"�y7�P�e�2B�F��kh�-b��3`���]�P[��
u�����O~ɟ%�ΣD�;�O�B VB�õ�o���o��l�Sܑ�j(�7H�����g�~sȊT���FrB���o�G����=dAE�Q��a�e?���X)�/0�::�T3<c�.�Z
��C�Lj���k�9�ar8݅�����O�/g�
<n&��*���Y���H2#{�!���#*�z���s�S�yMC"�e��:�yr���w�<.�X�(��M�s;�%v;�M��qN��40խ��t+��#�{�:��I�͌xX�ǂ�i�#L>�hL�vƄh��r+JY�����x�������$s��Cw#����Q��Fg����ɻKk)�J�w�Fl�B���=7"���(����J���/J�״�C��</�_"K�-�9���x�V�J��T�ȖO$�<�N2h�u/|��~�&���7 ��z�_K��L����r2w��>�Y�ޏp4��B߾=j�p�V�r�qZ���iΟ!ב������|��υ�j3,�O�\��,�z�b�C7+���>�����J����@���[��&͘Ne�*w=�@/�&���ڮ�߬d>1���pƏ�s��hl�v�ƎIÍ�<9sg�>�_N�1v������vȅ"%N��q�pl}^�,dZ���`C�Y{�${Z-�6o���ܱ 7����&���Y�p���~����L��#��e
��a�S�L�:��3���ߊ��V�<��P?�:�)()cvA�1kg�щ��s$`��4a�9`�'h^��o� �&���t�N>I�8�� �I�PQh�qgWOF�����X�����3��[�%G��z|~[Rό2�v�7;.�QɁT����e��0��M��0d���W�U$��5��Py��f�]e*���ŪY5ʸ�K�dOQ(.	-�o�w�5�%��L����3�J����a��Z����(o-�鿳)��l�5gBpC�YƢ����$x΁.���	{6 f-P�D|u���|�`ͯ�r�颯�'��3u��QV��֑P�{�7�#,�;��{�;0�'�J�J�H���M����	��dzk.�hK��2)jӭ��� �� s'BU�`�W;8Z�~�!�b�x�l�ATS6��mdi�ٔ[lk���/ƚh�Y2V}�L�h�v1�Mr�TM��t�h���'U��|�)�`w��4��;J&x�ѫ[_��}�`��{Ų����$fr~Q<��̸�����8q2�t f9�ȸf��R�y��:�u9��;�zl�4�5�=G�fP��>{goA�Pӄ���n#s>������κ�i$iK�f)em��s�ŧ�Y5�Of;���9�̘
���5��<;(;��o23{.���]%�M�u�LT|D/R������Mi8.0�KJ�8I6!�		�]f���τ���j9po��8,����V��yG�H�˧�#Q��r��䱽Ӗ}N�[lG��(ÀO���S�����b�=مײ��i����y�$9t�H_��t+Z�����F��3ѪvApm�~�2	@'�?#�����^g�ِ\"��w`2�H ����qgK���ӣ$����b�傡fr'��_�Z^V���%A_��U�)3ɾIt�Bxf�:!�Bs*}�����E4�m|�� �Q�!�d>M��p�`�^��:��>��gC�f3�DL�'M�tS��85:<s/	��>o�|��mKʈ�R�Iq#�dFg��#�Q����<����w�T�>sݯR*�<J=��aE�[�X��W���F��׍KF�/�9��h�Wo��Y�M�ˤur�ɺmh�=�G���d(/b�a��/J��U��I�q�/;ě4w�G��K�����3H.� =���ə��**[0�`V�|lq�H�^�r��Q�������#H��|����������l�W��f��.&eͭ`A@�Ľ-�8x%����ݵ}�܁��3�>wѵ�TF����`|&t��\xlO�E����l��E?���a%�zP{=Ā�Z��98�u���ka� �OT1C�ZhX����C��'�����]~a�)Q��6�����+�Ft1��@&<��M���~�?^�I0�?7.�~Pt�P���ّ@�D�oڧ���J�����FL�6:�o�,���_�O���R;�9҈��${��w=� ��{R;�'�� �8���'ua�p+Sդ�D����O[p��p�n� ��H`�.��YK�@[(i�[�[�e)oP��}j:{2��=2̧����:�����ғ�;��$�ɢ£!U"��j�&(qa�;�f�q8��Î�R�M�.�%0I��>�#������H߻��i\��\@�q J�&���\���[x�0��#��j��3�{Gaӏx+-�S6�Bwo��^"OM]�>�؂��E	P�,!���ؿ�{h��C��U4�'��B�H��&���>�~mU��UN�/�}�;�<����=m��4�]��DW�,�����e�u�V�f��l���]�v;�k�NGɻ�廙r�v�����T{��{^q߄.�2�W{#E�uen���qZ�M�uy�� �9���QQ�pR���¿J��	�B�6�b���~�k����$��֩zE�S�Ĕ���e�K��,K<�HN��
XP��Ü��D�9Q	1ߎ�W��(���H�.8�U_G^}�/h���:*Kr׊����n6�}��z�Pc�k[��y���ʊq��Kx�P\qAˁnK�6w4�L��a+��?u��gpX���B��]�L0�#�V�kNDYT�"6�%a\�X�t�rt�!�� �VdZ���\��5b�y�n����b�"��	n��ȥgS@�?ł-}87��x�]sG��M�1g��#E��~����	(d���^��(C��L�17Z���2LZ:����h}N�9������Tp[ �m�����&��&ݣeK�O�R�	҃��,�8G��5���8���z0r)��m�h4�@��줱E�O�ą1���tY7����2��
��m1:�&��1[��tx3$��r������Ps����n�Y~�Ϥ���>�H�k���8\h�~wD��y����58jH٤�ɋ��	����N�݄� �bkm����X��)e�w')c�o@X�O���� ���� ��Y�x�I�S�|��Ղ�4��e�$0� n����
���8��j��������ɉgR=��UK�$4���ڇ��Z�ޑ�%���%c�m�v��d�~�]�ۚ�QiA��M[��)�o �UH��cZԻ(�ѐ�{,[�X]/�&��:�O�5RӧY� w0ܴQ�?	C��ŕJf<��H�I�@�\W9-]��>}53��,��j�4�yJ��K�|}Yl'Ca��p� qk*����2R#�����7�M�7�ȥi�Co�� �DP/�����k�ˆ�{)��#"п�������2�ߋ�@��wv[k{�6G{�̔�]��M[mLB3��y!V�����t�h�B��_2@�&�`GhJT#������ 0?��Qި ���s���!���$����;�;5�+��pǅ �bn�f��ñu�i `�z����!f'� M�;�*�7���@�:WZ-Ļ���t ��)\������]� �]d^ ��X>�f`�I��Sm���1�(;���t�KfЬ$�`#7%>�,p�Jv Z)k�LCz����2�ŅyTN�C�nR�!v6v�JӨ�r������w�:��4Y�.�����Slb=����]]�ySǠ�$j����9�p
(�dR|��;��^Mj8X۲�-�Ӌ=���P1˗� �'1��-�TDl0����؟�U�y�}�}�}��%��3�8�/N�J�҆Xc5@ʇM�-������g�Uҹ��]���%+������gk�sTOJ�H2��uy�t���"!CJl�vt���W�����+�3��jG��J8��dK�7 =,QGm�0��ǿ�.i�(�.��o����� �$�J��2e�X#�lmv��#�Գ��C&d�K����Ae�⍞a��#߲�ԥ�+g��Hm�* ����A��!Ƈ�5�Z�I���KV)�-�>ۺ(�IV�B2[8��p���h�P=�#����r29i:7#8Ku���t%�cUV�^����R=�	(�[�\�N�]���H h��}=I��`�����k�}�N����'�����hT㦘ݾv�M�^A:ؗR����kg�dt�y�̥���c�*��2y����x��@��n�
���QL���v��%i���2�mj�Y~���E�<wͻ)��	Y-�h���Wv�ߵ�G�TE]�d(4�z׫���+������í-�2Ŝ�o�x��$�+[�勠Z)�QV�MC;��B�.�~F0��A;'
t@k�]�:���SI���:�'��|:C��b���(�R������<#�!!����;R��Cz��gV�G����wIfTs@�f�&�`����Z����5�&�a",�Sg0�ә!��^����Q����#�pE��V ��6����(�xz2�����6�ѳ}m:5�Z��P�m|H(}103�n
R�T�c,��~D�G�6a�E9g�p�;_�̵	u9��Ck��E�e���3�A	�%j�`�8�kp@��M	����U�r�����&(�D+1煞l�̌p��������?�{+��DRy�^�͌�c��wC+��bz0�s�j� T��U���n���!q/��$��<����?�������[�9R��m�f��k�z��.>��Ι��֔jiDYl��2x
�A��Y��.��i���2�-�S�݆��Z-4_�?�9�3�T{�j�9;ů��L�t�Ȑ!��Ud�@��.�X)�R�����+.r�	?�."� }��~R{jn��9ٿ�$6GiIuF�4K*����Ie�H�F��#�bF0�	Զקbx�p�'ܚ;S�1i����)����5��I����ٯ
�o�[��\�d���{�J,�޵����󡣷��D��V�x���Ղ��`9g��Y��N6[�6��S��	l����l�:E�|~T�V�����șۡ�������rԋ�8wa�ș���L�G8�:�T��I��5���*�2 tU�jrxĩ�r�U�,W��� 2�M;杸q:�n�[t���|��$ɬ����Ʌ%�"��ý����W�u���OB@x�C�A�S��G��S5�O�����ǖ���v9%����[��ֆd����%!4X+(���試�bx[*�C��wg��?~o&�$�h�ƛ�'��9�t��XQo0HC��9R�⤠����~¯�O�c��n�Xr��x:�H^�a`~��VS��5c��)����S	v��\�md��u8��q�ih�TL��d� o�;�=[��SC���7Es�{��`�.+h��+!����Ku�'�_�+��m��`ٽ�jwɉ$~3^�{7�:<�(����c�;g���J�M=Rg����z�(L�����{\�@O�Eڝ� �(�q$��,��O<4\R�e�ېX\y�I ��*z�\T����mkt��y/Q�����d��=�m̶<<.�x�os�/��o�~|@����.�ft�7��ET�3D���k���;2lX�oa�
:s�00@W�%80��&��w��j�|.��),`�P���j�ŭ������BD��.EB8��dm9�F�x���1��&<��B��2�)�"����[������nB�Ͼ�:�{���C�l�0���!�޿{V�:��/ct���䞟��l�ҹqpU���ҫ��� �kq�:�^TvBj��9s��s�σ3u
-�x���*K�M��c��@���Y�Xm:ف �Q&Q��ݺ)]$8@��������Ge&P��''��720k��j�D�h�Q)�Jx�Н��x\��IE ��V�G�m�^�u�$�cq<,kFiDͺ��9�u�upSu>3��	�w�˵��]t������*��;�-ƎRNRP���(�&i[<�#+h����E�4��͕n�+Ա,\ x�9�.�|�Yi�N~f�F�c�V�6�M#�73�"�$�+"�U7T?7����������8�r)���C��ˎxv|�[��]aVȱ�k����,O�;�smk������\)���|�uЇmv�)����1�^כ���v�cz���d��|��@H��wm�S=#Y���2 ��Yct�#�^95��~�*k�)�ܷ77��y��?up�Y�����K�������j[L�F�34�pmdR����j���Y����m�&���c2�r��.Ɉ7��@6%��<���-OoZ%���M2G5^]i�[�r��>&�1����3��� �k�0�=,o8nد�דO��Ŏ=��5��f�s�~�F�B�5���
�B;;���ܜ��%k�+�N�s��,rTJ<�!�%����G�����*�s�U������c�
���n�s%�8�U�&]K��a�&TdO�6UV鄗�U;\�Y���R����t�:*�6��*��!�Y�j�euD�y��L������ke��h�1��	�}�����{�C��"�G��3_F��0FP��5]�±b7�܀�&i�9,P�:f����zJz#�\�'M�u��̭~eZ���63�Pp�PD�D]|#>���S8�񔬋��M�m#ሞ�w���志�.N�lCW8@@iwf���O�l�{�J����vH7!<��QׅEIh��Y��_��U׍M��"�L��}E(���X��86aQ^�����w7�B�vW�FK?�������/Wg��?i�Yϻpx�)�#Ͽ8�*���O'�M���J�����6I�!��1=�c4c�~4Ns��o5��N�<B40	�c�����A<~E���_4iW�E]�<7eI3*{�u�(3F�' *�C�C��ι�x*�$xS-�e�
l��+Է˿G݆Q�l 2.�K����3Dh��;��y��_��?v��sK��\&��}�30se�-(p�?ٝ����ɒ(�hUt9����81J�Y��(1P�dO �a�t����gr_����!��g�H�S�tv�4V��,���M�r�~{�3�����ʵ$}.��ݱ�`�x����(j|�I�h[ʬ��s�MWBN˸���	��,���Nq�f�,�\+V���|�`T*vCbW����KZh>���U�ܟ��<��@�Įtt�!��{�������TGa��o��r���ʋG��M.�d	�0�HN�^�~�;����]#��.�|�{�`�yp}��0^�����G~.r�XZx��jt�k,`[�|d�b���o�1�IpV�O(Dx�E���e���F�뎠1�䳬��T-B�M\�r�泈�c�Jș;��:�[kڝׁı`�oi�5S���8��YSck罹@����Ȓ3RCD {k_,�����N��0����>h���[���G�)R�f�ٖ7˅�S?�A����]U�7j�%��G�g7������6��&Po����V@�X>�����1�}�ur�ÒE=�2K4���2#��y9�ox"��o�Y�לN�'#��3����ri��~=�2�2T�$�6�����F�����\�r&cϭ�э&)͋���JE�l������.�T�����\�S������4����U����I�mz������Y��V�t��s�I^�8A�����	u���ǲ~��cF��U��m���~L��A���>�b��6�C��ѡbT�̽��_T��� d��ֆ��l�L͸а�K�����{�9A,^�Y��h,��"X_V6X�ֈ����r|n�_����p��;Ӽ5�AUI<�O��Z��a�|h��\�qf�Q;�G}M�Maj�f}�I�{���S��A�.cm6>=���g[?N�W�֟紫�����r��>_	D��xb�������ǀ��O"�G��J�\���WJ5��歙�Ä/��H%�S[�Z�a?��:��~���:�- �Vq��kCI��6{��������w;�1I��>�7g�T���4����5�����9��aw�Y�Ц����][u
 �]߀�|�t.^��a��}O��ɣ����S�4z8l����g�+V{n	���kQ�o� r���؁�>���ݣ�z���v�Km?��~�w5���|��R�
17
2�
L�P[�T���������{�5)�|�Τ�����=)�r �0�MFS�p) C
����9��}6�hH�l��ovhz�8;�Y�+Rec����ѬQN:�����R�+�_��.ǰț��텢�K�(�J���O[_�m?'QS�ǅ��%P����<�|dp�O�� ��� [IR��:��G�����w�x[���Ԝ��j�T�-�zg���E}x����֤����B~��}[d,x�hRB ���������co�oEL�5��������م�� ��p���Q��&�>����z��z �w�6I��	�;�P��:X�9)�͂o/���_4K�9�N���t�U��UƧ}����7
�_�M�^���ˢ�8b)��+�4�6Pq.���2�����4��AU7v(�2�+��hI���\�����`*��A�]�|5	L]"�_�����V�h0J�y�9i����5nk�|��mK����gA[����dMRH�w�sr�=�)��ux��6+�Rs'��6�-��:�>�o�u&p̦�>����[ҷ'vA��׻���c���{����EsK��Vb+R!�);�J����<�Z��tvG>ͭ�+`,݉0�M�r���$���W�$���(G0��$F���Y��C�XG7��� 91]�9yS����:�����N?�`��r7z(T$��iQ�v��X&�/lHŕ�0�{$�˒���x�
�o�:�3<����{���c1Ȃ#(q�u�b�b�C�Z��Frg����t�6�����ڟg���|W�}zU����P��HL��9s�	a�լu9ZnP�Ŷ��
�U�Vb6�bC5� ��W�mƟ�aB�>����E�j��<�H �Q��c�$�?���>���j�(*��~�z�@l�&I
0	��{��/�2����rr�2no��S��E���#�э���[�.n�B�W���\j�^N�*�J�r��9,�ݦkW�$&!�3�#Y�Eű~�I�&kc�:�L�+/X��LL'(�����$I�G�"��[_��:�����J8�T����di]�kpM�&QV7��(�<�c�8�V�atb�@���c�!������X�A�[��(�$�wƋ�1�E��Ȝot2���O;~.��	9�:��b��Ԝ=����V�����K�4O(������(��ݪۙ���Þ":������iw�"?p�L�'WJM�f`�SEyڤw�A'-�ΐ�,��U��֌3yp=+��C� �=��y���\\����5!��Fs�3h��̍�q�q!t�B�`S�E���z�p�&�.�"H���tt���D4|+�E�@b�R��{�뻔fY�Y߂��[�����+�!��/��>�����v��/Ww�������}���X2��39bZ$��z*bg��N�U��� k*2��H�S�uY���[*ʞZ�"���|�xd�q
���'�%��-5�d�,�:�`$� >��|���M]�1�h^����ܮ�ݼ� f���椄�:�&�����rFc��hg7��ɠ��}��6=����5)?��A��)�'�G $`J��޴��蒶��i � �����X[J�Һ$�[~�I�_M���X!Q<�����=M"����p��2l�bB�a�����d{#�@���f���\�H1 �F�-(@.�ڝ�IE��\�ѣ~�� uVE*eS��, Bck�N��p�K���P�G��?<en��/ӑ������_Y�q�R��=og�RZ�)��	=�.��،���̤��~NF�-�_����ȥ���G��i��d�؍8A�2�@�B��?d ��[�3̵zr�P"]T�,Tk��s�\6�Z�~^����[�l�@^������ufJم)ԕ����b62�riD��BȒ���A?�(�dw�9L���À�p���L ee�ަ�ME���'�����=%��}TZs�y�h��	�ӽ���i	+�UUu��(�O�./����~֣�L�C�H������m�����I�*��xc
���6Z�u>9L����o��'�^?���a�"=�0�,1]����cy�s��yk�Z�v�\���4� 'p�Ε�����BpG*�����Q�U��	�( �ԛ�OM�Z(�vm�rv�VC���k*O���b-MC�!]�r�.q�S'1��TN&���i�&�jy�5,�y�#W��ę���a-$����+Neȥ�j���f�	4�h=�,�1�ůQ��"�@�n��܎Fi��~b��D|��J��aSwK��ZnG�S���p��E��W��]]27��I���uMr��o��yd���UL����v��O^����ؾ��2�І^�'f��ѡ 2^�~�b#��нA������(�\���©��XY�B	(k��{WF�Ė��ɕ���*�zga ^���
_����O8���W�K��n�W��$-�_I�=,�����3�"Z,M5N0Y�UW��Ǒ���0	�B�//�*hQm��׈Ca���<�BCx*<@qNK4|�����l>r��G,�mT9z<{��[} ���4{v�z��EV29講��m��W���V%rC���v�v��@m'��K8D���[�n}��3��~�0�&x�3�C&A�V&˥N5���y�!l��;�o�.�Y�I��7��Qʳ`���w��f�E�#C��y$�oH
o�hXO�p��mY?�T��T:1q�C�	�Y�������ϲ-x����y�����ѦsɏЎ_Ao�Rn��)m
[mB�'�7� ��?��R�#G��u\c��v|?�:6��6��[Gկ�;��gq|T���[�H��Z�!����H�Ս�2O���%�'9�sƩd����N8����w���ic�/ш��}w�c�<`�'2-Ĕ��V��Ll���Y8�G�V2F<z2
8���y��B`�maSC�z"�;A0�^;<�xz�}H��Ⱦ��s�s�s,
��g�B��rğ?� b�8o@W�8�
���"�Hvs��n� �7Q�"�fkɷL�G�����c"�e�s������,���OT������T��"��)ed,3��β��u�/���DCH"�S7� Q����������Q�|���=j��v���Gly�L����Q"�ľ���41Kp������BFoz��\Le�h��B�ԑ�0�� �nF���J�&�J��$��Pb ��e�������>.f<����RF�g�3��� ��q9�#��̈́�R���^q=�v���oZ7����a�?��?�g���e-�ޏo�1�N?A��6��e�s�>tm+7��k��z�����	��4�Y�\�]����K/�s�=�L&����{?��Z�f:%*��⡝���� �M�=1lZn�C� ��3��3G���~�h-�t�d�gY6����,?{V��}���E�F���+b�l����Dt�� &)����M��*�j���`��������mǄkA޽�e4�h�NTk[�g\,�8��	��i).�웇J�0��ϱt��wO��Y�Qù�(p��`�]҉1*R'��XD��F�Z�ڢw@�+�S��>�z��U��;x���]U��Ӧ.2ܨZ�ų<��*�Q���K��/� ��	��J8EZ�'+9�� �5�tw�F�e�~z�:��m������(�!�\��ތ���3G��������kA���0�f>B4�O��Y�
(�T�`��ߖ��wQ^[Ȃ3�A#em�6�=����B1I��e~�f7�0�6 ���[xL��Zp:�y�Ys�R>nJ�t,�@afo�
|_�u ϫ<��]���,�:���e��Q��#��=A,���@Cy��[������Zy�;���R��ؑ�H:`<i-�LN�)j~�pp`/�2���X�WY0���1\�;������.��d������E�i�^�WkY�_x`�'�v{�m,1�QP��[u�	v�QJ���=d�� ��<�����|���m7D~H��g#&1B,�GiE�W,��i"�%��dM�Mh�0ޢ����_ԁ~�(���CJf��, �M�ێ��D-gp$�or�!NW%fR��=���FƩ���cMy�Y�������4?xp�s+��`�3���.eS*�?n��P�PwJ�`��^��ʱ����)�C�� 3Z�#��ȹB��*�Q��d���G�W�pq؛��!���M�(g���ҭQ�W����:Z^�%티�o��e�AU�v���7�Z��e����9��(K��B[ߩ�E�$�t�+����|%�!����Bp��4�H�	�t�5�?,S9�m�%R���>�z��=5�?:��r;�LWed�����=R�
�<,:5�VA�u�6nFYº��Y
xٖ8Z�m+��KW���Ymz�AUQett2��u��yQD��\S�������eƣq3Pm�r�2k��@����4�ХI�mI��p�&��
98���j2��fJ-/&DD�U�j�\�b���N��h�av`oz�"(F��:�Hb�n?��/m����� !k�1n�n7۹ا�{r#�='.��n)ݿ�a����gZ̋HK+`<�>w�&7�t�S��3W�EB�x�e�=����ԣ�8H1�t��NFa�1�ˎU�G�������zpn�����S�Wkj���~r1�s��H�A�a�NLIŔ����o�΍�,���}:ҹ����~x)P�]q͹��d���K�6��3�8���ӱ3����$\��h��_[};9�c�x[��DXȴ��4�z��QV��i�شG����jD �?��QY�9'W��ETT�ɉ�Y!�x�My���l1#�P[��qe� �����N�q��3y���1j�f.8Bޞg�������
�TF�r�S�Z���x}i�~��^?���_��3�f�Vs(��hV~���V{��� ��x��*w	J7�ܹj>�g��X5��;��x���@dw��=k�K|�5�����w	����T�š�c���j�й� ��a������\ɗ���#�N��&��}-����@��^z�X۹=�ܒ&�H;I�*+ha�O)�t��ٺG�-�E�!ZR�Z�B4�{����<�ہ��/Z��*�L�<�y��(1��:l�,-ˇSv��oG�'A����ZB{�83ƈI�-ԌXl3<��������A��(�x�Z�:P���n� �h�zRWGfd8�\�椰�Z¹2	�tΩ����_:q(�3���ܲ�QRT�%򡿀�"�L�V�I�������������)ds#�k��C%?ż�
f�4i�����`B��e''m7�΀�2� =��u׫��*�1Ѡ��18�'���ECmu˓Е@+�����C9�4+����BH$F�a�0��O�TlW���za.b�0_>��Ʋ��Q���87�
Y N��r���`9v[D U���^7���v˹x%kW�~��hD��҄��k���k��ꏄ�3�1A����og�+[��9��'��
��2����a��Q�g}"�����k���|}��m��avt�Ɯ�Iիdq�j��,�w�8�.L�r�A�<χq�W(��=:X�?��������I͠ϗ��M��)c�	�1��\e�S��}��l$���B�"�Jc(&8��p\��?Q�e��S'�F��q����P���~I�I*-v�Yd�I ِ��n&&'�錑�S��vf��VB萝�RJn�!`��h&�9�� m[���T79ã�h����	���F�*n�T�"��iu�J�0 ��L^��ӗ��.\	�:͹�t*�z������xZ�f��b�)9V���]꫰Rٳ�
 ��t���:������{v��&����� j�	1�"N$MZ�ʪ���K�ua���>>�<J�d'*�Hr���ҏљc�c9K���^�W �3�<�#���Uo�����dr�!�?�:���I�754W���7�|T�z�������:�Q��K|��JY�%PE�Ot��Q�O��!̬���ץ_wao��g�?&������Vj{�B���_����7�j�uU��H��`��Y�GK5���2�9Ԃ��Y���K��{�>6P~�Bй��D��,#vir�*<�ۦ�� �**�V+���H�@�:=�x
��n+S��.����w"�L(��;�.}��z��swg��#�N�M߫46l��st+���KT���b��Ƌ�h����|����{��c0�K���>��Fa���=B^ѽ
OAҞ����t�-�?��p`~<�#�d�cgEf���Q`3!�Ԃ(�u��ݳu�U�-7����+�v�z�U\� ���4��!#�H���ZN����n�|�D�kb�ת��~\/j�47k�x�4�Z@��Hh�'�e��س��WB�Z)����
�2����>�e�'g�Ĭ�@�@��SG�Ŷk����tkb�;�h;^�ԕ��v��ϲF@�u����!Ɔ�o��8��Ѻw���	�:��޿����fu�~0��(Qdv8~���������H	��1��~ؙ�C1|�x63�g7�wZ?��>E2�
o�n�RD�`����3-]v畛h�o0R�:wm{�6q�`�CI3�70��烆�Q~x�K"E��/}���2H��MS!��wwƆzß3{M�k�˹�!H��I�����TD���}��-xx���"bWB_��BR�B��]�W�쑂S8?!X�f�tkB�b��᳹����.g�f[�6h�m�v~��O�_�`<7|�b�r��s*��N�����.�6]G���f�K�|����iظgۋ��$aڻ�ә��Q)G����EO�N��:�$XQ/Q*v�f��|��#�?ԽVJ�[����Ǆ2�U���x�ԆuD�1壖I`�-�73	�y�i \I�6̟�&_TB��vC���3]��xlnԉ�kp�@��j���5+r/`(k������<<"��y)�=)�-{������~�~u���(O1LO���'�Ds�����;0��im�rJ,��o�'�}>����)>?g�m�옚(����^G����Q�[5ȩh�緥U����&Z���`gu��b�=S�����֧0�ܑ����p���P�U:���{�9#�Zs�d+�������Eӂ_�=/��"b����ӿU���e���^�6�@�*�,�vCM2�Y.���q�r5����/gQJn���>�� +�?'Ql�+��9��r~[�c�AZ\]|cP��3s���CD]wW�5�dg{�K(�[N����^��8�V<�KN<��M�m��4�9>5�~A�c�ӟt���I�R{=���)a@0Q,|�����34�r���"��xf��Ù�\O��wR�'�q=`�(��w\�C*���.uH�PȽ�wM���܊�_���|�7�V�`��������Y [K`��ͲKD�eL_Jܭ�vw���I�L��}-4z��:���y���җ�H��/�Ph�wK��A�-vԆ��>�?���v�|��r�l�q]��rs��5O|�^���~�T�6��K���뵧,W��vA���"[��ͧke3��t��-M~�}�-MD8x��(s��$N}��'��������9L���&��Z�dQ9�e�\���$���2jD_�*4�t5:5-�a�x�~h�N��9�氾�g��A�����GR��_��@x��Ѷ�!��e����G
|(�*�Ri��L��� ���W��9i}LH��{p��9ſ��i��;Zb�8�� �$�X���r�フE$�5�c�kG�K�-���b-;0q��ザ[���!Av�h�vE�N���|l�e�P�y�H�Qc��8�"ɭD��j��p��6wQqՖq�N���'��G��j�߈l���6.J�`%0�;��ɼy���<�몞ok�(Z�?��E��!��F׵9������.t~	��Ml�� z|:VO"'@ºs#�i��'�ET*聎s�Ҩ@�.i�ȼ�^5�Ӎ9�7��Z�
���G_V!Kph�=/1�ٺIY/;�^��z��n�&��C��κfMh���8��A���?j%��m��U��oA[*v����,�����n�m�v�"�Cy�рH�K�<�N�t-�O<�_U.�����)y׌��X�
P��F`�uAj��Rw�1>�Ю��F���$�X�{�@���$ؠ!����\Gn��x�W����u M�6��K-I�(�^���0h4"�����݋�G9��x�ye,�G:�[<�Hyf�FCΡ�ٹ^�f�R[[l�0�:TY���rn�cq�� X�ȭ�������N���-OY�`5Q�>��ྠ��p�f��p��n���P�� �k��5�5�Y��Cl� �Re�d�m���;�兡�c�m�����f�jKw��v3��G�v�4*H��5�>ܱ��Nr�7�Is�bwń�N��.^~����l�=R��ꣅh�hhi��DG�f�0�p.k�?݇(��lۋ
�϶�����E�88�+� e{�W�r�f90'd"	�3����)zH����qrt�3��$��4�6@�� :�U61	(�n6ji�e6��.�1.��J?ջ���9���	^XB'Ї�Lf9��झ�uЧ��l}���3W��U\�!Z~ӗ��(�%�d���W��w�7�of�	)�����)^w���C�u�'_���Ol�8�E���(�?�����-f�!������������ywQ���~�1x3��In'�ލ��u
L
Q!j��#�"�4�Q;�"��*�g����R�z}m�(?�_�xN亝��o/8j�L���5�Ҿ݃�
��ѕ_��n��������Q.��l��K���f`B��Ň|�|�#?�/��6�a����0k�]�C Y��4�roT!^N$����ڥd�y&�&}A�㋡�$����E$�_bHL�t8�(4iq!J)�3z�&��Yp-n��m@�0������}��e؁	/�M �]y��;�_���0�Rq�]��RL�:�.!���)�՞����t[*�[�M5��v�����ҐѵŌq���yD>�4-F`���C�iYdz��>�ɹ��{� �-�9_��lr� �)�ѡ\:�VYwV����v˾H6��<��JQ/�&���q�t(�}ӛ!)&� ]�ƝK���Q|&s�r���S����#���%��"K��7�-O
��/�g�1=ĵpj"F]-�Q,�t��� ��C��'Z�|�$NE���?P��1�9�P�<z�����CG'@b��X�R[�oP�lNWm����:�K�㊯khr"��X�ܞ�1I��qy�!�{wX�ybyf���=|��ķj($&�+�0�A��@B�V���]����Kr� ��3�=��MF�lv˷��j3{,V�.��8�� b�43N�%�uF�Xe�SGD5��V΄H/�g�㭍ޯ⭓��e�8��� ���f�w�
��/.d��v��h9DƐ�MS�[JL��f����SЃת�t�ͨ���I9��#�����4��>6q���k" 7���ι�I�ã�	46y52<h�]���)����m�ۆ ��U[:RR9/��#��<����Y.^�� �
B��{�J�S*���*"�]}�ѣ*z��D����:!��Giy&A
��������HL��ݷ&��TT�ҹp#��9ĥc�AҨ*��v���ץ�A+��/�o�ﷱZRم��s�����j*R�)�:.e�)c$Ff�w � �|0+M>"��U��c���L�1�R��Q�j��>�69��$�B�VJlśV"��G�)+ښ ����ŹYFQl}��,H~��<�<�a�we�`),}U�H�=8V��h(�B�:u�q�A�ƿ���;3J��-zLߵ���8H_�9���� �vA�t|�E�$# ���W��!�-�3�Y��o b2#�2�=�t��4u��+��;A��e�|L�Z�7]M�֯v��~�w��!�Nv�D�Y�t�y2�δ��g
w�^�?O=��,X��8rњ����r���g�x2گKhXx2�#����!�>ǽ������kstu���/�މj"5��Nok&��M�47tߊtɗ����O,�`=�E��5��v5��1����+�7��W��VL�kL���E
?|Q�fɑ�������W����>���2Z�ǩ�"�fOY?� �/P��l2aѬo�A�k Ŵ�k?g/����&g�[f	�PU��c�>�8tQi��4䝬�0��ŏCد"j���n��g�Ҹ��N1���j�& �{N�S�A�5Y��'�`St�!��߽E���8{�q���2�h���ا��A�\�'�94�Ƒ��p�jl�{OzV</äY��gy(}O�V\�ąD�P�鐅����Lmn.�
�P���e�v-��A0�Fŀ{qy/C8�ǢO���9�
 )_��YGom0����s�d 9�tkl��cǛD ���?�{O�]��Oc���+a�� ?k!1jo���=�#!��3_*�@�*k��v��Nc��F2gm��e���\!*g�,�Og�kRU������������A��=L�y�]aY�=�L�0k<� �2\��rgL=���`%4qٯ�����i-a�����1S��W��p�Ax#�_¿��r�%�.l;V�ا��op�+��?���U���\.r�{��2͟I���_��mSr)`i�������^kp��x�q�@���$��H�=]�8�-iP`iP?Fy���ϡ"jGL���F#�[�D�Vg��v����H�i�L��b܁����LNc�V�ݖӖg�Q�f���e������c����+�j�+����*9�:iJ���\d~�&aP�������`�^E�;�5rݐd��   �A�h	ܫ$���_6�l!�$}hè@պh��>$�WV� ��V �RRlK6*�y���K'�R�����`Y��1ʢ�~�d6a���ŕ�rF:�ս��(㔰8��ݯ��Sʥ�\�N)���������+�ޒ�^�����8�ӃH�2J��o��b͎;R�~r(X�Ϭf�n�[�=�n��"��x�O��G
��8�aػ�"{�U<���Nm4j�p�ێy,F�1�G���0k�=
�P}���� b�̭8�����θ�y2z����]��M1e�Q�� B
���(pf�GH �tb�e�Ar��%u������z�f��4 D:�&긚25�fg�(����ֵ�mCP��|���mr�N�h����(������ĸ����X�E��`ݚ��*t���(fn]^�{�Zn�`�_Û�B�Y:�E͛�1�AX2�T�)��o��
I��p�L�����C!8�f��~�z�3�"/^ӡ�
Uj�S�,��o���� �ˉ-#�#N����w��\��[8�fBM���$ׅ���ZtSPZ�#s�.�������:��)$aȳ�y�����C�s�	d������a�'^w�%���pꤸy�? _2��<��'��(�K5�>�>�Xx��a��rJ�y�Xe�Jj(���m7X n�����ej����O��A3J΄X k��KG��W���D���韫 d�^�Hw�0JX���pkVZ�@h��,��(m���d����}�#��_)U�,��6 �y�C���}ˢ��h�WD`59�U�����e�r�v�-�I2O3���X�{D��$��aw��ڑudt�9����ڤ徳&��Ek�Z��L4���#ᩳ'�L�a̬�^5�]�<{�e���~���B�+JӉ���`�����9�,�)�`X��CNL��8��e@ocX�mU.Qt�����Kn�����|�(r�wّ8��0���+�^w���fS��~��ʳU&�E�H�K_�5]�P��ŨQ���~��o�Z�qG��@x��S�&�[4��A�}�(�u`�#�,������{����=Np>�����7���H;xv�.K�g�m������M�.p�'ȯZ.��0�%��>�E����a��&;AL3�L���5��5Z�T��9>���t7�I���lWsa�{��
,�o8�zu�ޱ������Z��_��_�ja��E8�v ��M�mg�R`���6��8��F4��oDz��:���&2�=�!���H�8��,$�il��Y�gw�C�L��5��Y�U��(�J�Ɯ,�.`^�!6B�e�ڊK5{�*͈۹�W���n�b���Y�E����f^��r����{�.�3����YT7��>�ps�p�z&\���+�-�j�}p�T���'Am�f����e&���g�F��UKM��T�����ɇ�>��l���XB�M�;��{u��G�{u��K�:}�%OY㺜H}����tra�f�k�%~�	�%��]=V��+�?Z��.S	�F��Y!+E�E	��]������}�{�P�fͯ2m�ǭA��#r`����ݻk�[R�J�ADņ���|WE�l,$4�@���x�&U8�s�R��GS��%a�㺢~��)�$"͘�F���x&����;����Q�@0���\�p���h!��U:�-�	2h���O��w���L�f?T�Ԇ�1���"���E�9�
[C{�
G}$BlD����������,y��ҕ%�r �*�N�3׍5�g9�����Í��Dm�Q0:��}� ��f��k�m��5���Q�e!	p��J+�m�v�H�ODy_&��/;Z�����MYg��?��N!#W�,B�ۣ֏����q�\?#)]P�hW�r�/�AuR�xSQ���5�,^hlBPt� F	�Cp��t�l2z��h��E�����k!>���b�'��=��æ�Eq��R3���t��@��J�fC�Nt�܋c��dBP.�\�jA�k���E�U����Y.%�b�l�}Xș��,,VE���`)f�5��j��v�����͜�m~oU�ixG@���
��|eGV|s�Z ��.�������v$����/�U�ꎄ�P/WΩt��ݨ3�Qԩ�hz�W�{�a�����	���~d���k�,q@U��#r~����&�����������iM6�&��I��H����vh�@��-x�Ո��zk�Q�[~�̮[������G�ݼu�Q�� �s��M��7��:@!9dDf��G�����c%��q����WTFB 2!`h�q3��kT
��9�(u��3�n@�'����Lg��j�v�Wy{��L���H�",-"���=��:��:2�����	����\�Y����r�H����Ӊb6궮�bZ�%��#��NY�C�y��e�l�������l+7>/G,*%�\�([
 �M�Au��V����&D烬�lN��6��u�#[����ZL^��-��!Ē��� �u��ѯ'Q��erN�*/�KP�Xc�*��'ڃ[���X8kO�]�,ҿ.�SI����.5b%+]:����I�:��^p������ܡ���Y�#�uU�u/�FLI6�0�\�jY��46��[�$�(v��F�os��x>dk)��+�r.��)�7QK�5� ��wv�z�X�ܪ�7��_�W@���y�Ɏ�.�(���u�-i�
�X�����v7�tp�@�4��B�Ba�k2����4�hcn���[C��7~���i'�:�[��p�i���)���d�SZ�>�A�����|�	`/�S'�i2���MU,��)�[��(km�T�e��T ��Ô���#�����~���q���l��pE�D]I�R�>��°��L���/b$߾-Z�%�v9Ì�>ARAk�>�B5E���M���