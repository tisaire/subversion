// Nios1.v

// Generated using ACDS version 11.1sp2 259 at 2012.10.25.17:30:37

`timescale 1 ps / 1 ps
module Nios1 (
		output wire [17:0] pio_ledr_export,     //      pio_ledr.export
		output wire [1:0]  pio_dataread_export, //  pio_dataread.export
		input  wire [11:0] pio_data_export,     //      pio_data.export
		output wire [7:0]  pio_ledg_export,     //      pio_ledg.export
		input  wire [17:0] pio_sw_export,       //        pio_sw.export
		input  wire        uart_external_rxd,   // uart_external.rxd
		output wire        uart_external_txd,   //              .txd
		input  wire        pio_rdydata_export,  //   pio_rdydata.export
		inout  wire [7:0]  lcd_external_data,   //  lcd_external.data
		output wire        lcd_external_E,      //              .E
		output wire        lcd_external_RS,     //              .RS
		output wire        lcd_external_RW,     //              .RW
		input  wire        reset_reset_n,       //         reset.reset_n
		input  wire        clk_clk,             //           clk.clk
		input  wire [2:0]  pio_button_export    //    pio_button.export
	);

	wire         nios2_qsys_instruction_master_waitrequest;                                                         // nios2_qsys_instruction_master_translator:av_waitrequest -> nios2_qsys:i_waitrequest
	wire  [18:0] nios2_qsys_instruction_master_address;                                                             // nios2_qsys:i_address -> nios2_qsys_instruction_master_translator:av_address
	wire         nios2_qsys_instruction_master_read;                                                                // nios2_qsys:i_read -> nios2_qsys_instruction_master_translator:av_read
	wire  [31:0] nios2_qsys_instruction_master_readdata;                                                            // nios2_qsys_instruction_master_translator:av_readdata -> nios2_qsys:i_readdata
	wire         nios2_qsys_instruction_master_readdatavalid;                                                       // nios2_qsys_instruction_master_translator:av_readdatavalid -> nios2_qsys:i_readdatavalid
	wire         nios2_qsys_data_master_waitrequest;                                                                // nios2_qsys_data_master_translator:av_waitrequest -> nios2_qsys:d_waitrequest
	wire  [31:0] nios2_qsys_data_master_writedata;                                                                  // nios2_qsys:d_writedata -> nios2_qsys_data_master_translator:av_writedata
	wire  [18:0] nios2_qsys_data_master_address;                                                                    // nios2_qsys:d_address -> nios2_qsys_data_master_translator:av_address
	wire         nios2_qsys_data_master_write;                                                                      // nios2_qsys:d_write -> nios2_qsys_data_master_translator:av_write
	wire         nios2_qsys_data_master_read;                                                                       // nios2_qsys:d_read -> nios2_qsys_data_master_translator:av_read
	wire  [31:0] nios2_qsys_data_master_readdata;                                                                   // nios2_qsys_data_master_translator:av_readdata -> nios2_qsys:d_readdata
	wire         nios2_qsys_data_master_debugaccess;                                                                // nios2_qsys:jtag_debug_module_debugaccess_to_roms -> nios2_qsys_data_master_translator:av_debugaccess
	wire         nios2_qsys_data_master_readdatavalid;                                                              // nios2_qsys_data_master_translator:av_readdatavalid -> nios2_qsys:d_readdatavalid
	wire   [3:0] nios2_qsys_data_master_byteenable;                                                                 // nios2_qsys:d_byteenable -> nios2_qsys_data_master_translator:av_byteenable
	wire  [31:0] nios2_qsys_jtag_debug_module_translator_avalon_anti_slave_0_writedata;                             // nios2_qsys_jtag_debug_module_translator:av_writedata -> nios2_qsys:jtag_debug_module_writedata
	wire   [8:0] nios2_qsys_jtag_debug_module_translator_avalon_anti_slave_0_address;                               // nios2_qsys_jtag_debug_module_translator:av_address -> nios2_qsys:jtag_debug_module_address
	wire         nios2_qsys_jtag_debug_module_translator_avalon_anti_slave_0_chipselect;                            // nios2_qsys_jtag_debug_module_translator:av_chipselect -> nios2_qsys:jtag_debug_module_select
	wire         nios2_qsys_jtag_debug_module_translator_avalon_anti_slave_0_write;                                 // nios2_qsys_jtag_debug_module_translator:av_write -> nios2_qsys:jtag_debug_module_write
	wire  [31:0] nios2_qsys_jtag_debug_module_translator_avalon_anti_slave_0_readdata;                              // nios2_qsys:jtag_debug_module_readdata -> nios2_qsys_jtag_debug_module_translator:av_readdata
	wire         nios2_qsys_jtag_debug_module_translator_avalon_anti_slave_0_begintransfer;                         // nios2_qsys_jtag_debug_module_translator:av_begintransfer -> nios2_qsys:jtag_debug_module_begintransfer
	wire         nios2_qsys_jtag_debug_module_translator_avalon_anti_slave_0_debugaccess;                           // nios2_qsys_jtag_debug_module_translator:av_debugaccess -> nios2_qsys:jtag_debug_module_debugaccess
	wire   [3:0] nios2_qsys_jtag_debug_module_translator_avalon_anti_slave_0_byteenable;                            // nios2_qsys_jtag_debug_module_translator:av_byteenable -> nios2_qsys:jtag_debug_module_byteenable
	wire  [31:0] onchip_memory_s1_translator_avalon_anti_slave_0_writedata;                                         // onchip_memory_s1_translator:av_writedata -> onchip_memory:writedata
	wire  [14:0] onchip_memory_s1_translator_avalon_anti_slave_0_address;                                           // onchip_memory_s1_translator:av_address -> onchip_memory:address
	wire         onchip_memory_s1_translator_avalon_anti_slave_0_chipselect;                                        // onchip_memory_s1_translator:av_chipselect -> onchip_memory:chipselect
	wire         onchip_memory_s1_translator_avalon_anti_slave_0_clken;                                             // onchip_memory_s1_translator:av_clken -> onchip_memory:clken
	wire         onchip_memory_s1_translator_avalon_anti_slave_0_write;                                             // onchip_memory_s1_translator:av_write -> onchip_memory:write
	wire  [31:0] onchip_memory_s1_translator_avalon_anti_slave_0_readdata;                                          // onchip_memory:readdata -> onchip_memory_s1_translator:av_readdata
	wire   [3:0] onchip_memory_s1_translator_avalon_anti_slave_0_byteenable;                                        // onchip_memory_s1_translator:av_byteenable -> onchip_memory:byteenable
	wire         jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_waitrequest;                            // jtag_uart:av_waitrequest -> jtag_uart_avalon_jtag_slave_translator:av_waitrequest
	wire  [31:0] jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_writedata;                              // jtag_uart_avalon_jtag_slave_translator:av_writedata -> jtag_uart:av_writedata
	wire         jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_address;                                // jtag_uart_avalon_jtag_slave_translator:av_address -> jtag_uart:av_address
	wire         jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_chipselect;                             // jtag_uart_avalon_jtag_slave_translator:av_chipselect -> jtag_uart:av_chipselect
	wire         jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_write;                                  // jtag_uart_avalon_jtag_slave_translator:av_write -> jtag_uart:av_write_n
	wire         jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_read;                                   // jtag_uart_avalon_jtag_slave_translator:av_read -> jtag_uart:av_read_n
	wire  [31:0] jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_readdata;                               // jtag_uart:av_readdata -> jtag_uart_avalon_jtag_slave_translator:av_readdata
	wire         sysid_qsys_control_slave_translator_avalon_anti_slave_0_address;                                   // sysid_qsys_control_slave_translator:av_address -> sysid_qsys:address
	wire  [31:0] sysid_qsys_control_slave_translator_avalon_anti_slave_0_readdata;                                  // sysid_qsys:readdata -> sysid_qsys_control_slave_translator:av_readdata
	wire  [31:0] pio_ledg_s1_translator_avalon_anti_slave_0_writedata;                                              // pio_LEDG_s1_translator:av_writedata -> pio_LEDG:writedata
	wire   [2:0] pio_ledg_s1_translator_avalon_anti_slave_0_address;                                                // pio_LEDG_s1_translator:av_address -> pio_LEDG:address
	wire         pio_ledg_s1_translator_avalon_anti_slave_0_chipselect;                                             // pio_LEDG_s1_translator:av_chipselect -> pio_LEDG:chipselect
	wire         pio_ledg_s1_translator_avalon_anti_slave_0_write;                                                  // pio_LEDG_s1_translator:av_write -> pio_LEDG:write_n
	wire  [31:0] pio_ledg_s1_translator_avalon_anti_slave_0_readdata;                                               // pio_LEDG:readdata -> pio_LEDG_s1_translator:av_readdata
	wire  [31:0] pio_ledr_s1_translator_avalon_anti_slave_0_writedata;                                              // pio_LEDR_s1_translator:av_writedata -> pio_LEDR:writedata
	wire   [2:0] pio_ledr_s1_translator_avalon_anti_slave_0_address;                                                // pio_LEDR_s1_translator:av_address -> pio_LEDR:address
	wire         pio_ledr_s1_translator_avalon_anti_slave_0_chipselect;                                             // pio_LEDR_s1_translator:av_chipselect -> pio_LEDR:chipselect
	wire         pio_ledr_s1_translator_avalon_anti_slave_0_write;                                                  // pio_LEDR_s1_translator:av_write -> pio_LEDR:write_n
	wire  [31:0] pio_ledr_s1_translator_avalon_anti_slave_0_readdata;                                               // pio_LEDR:readdata -> pio_LEDR_s1_translator:av_readdata
	wire   [1:0] pio_sw_s1_translator_avalon_anti_slave_0_address;                                                  // pio_SW_s1_translator:av_address -> pio_SW:address
	wire  [31:0] pio_sw_s1_translator_avalon_anti_slave_0_readdata;                                                 // pio_SW:readdata -> pio_SW_s1_translator:av_readdata
	wire  [31:0] pio_button_s1_translator_avalon_anti_slave_0_writedata;                                            // pio_Button_s1_translator:av_writedata -> pio_Button:writedata
	wire   [1:0] pio_button_s1_translator_avalon_anti_slave_0_address;                                              // pio_Button_s1_translator:av_address -> pio_Button:address
	wire         pio_button_s1_translator_avalon_anti_slave_0_chipselect;                                           // pio_Button_s1_translator:av_chipselect -> pio_Button:chipselect
	wire         pio_button_s1_translator_avalon_anti_slave_0_write;                                                // pio_Button_s1_translator:av_write -> pio_Button:write_n
	wire  [31:0] pio_button_s1_translator_avalon_anti_slave_0_readdata;                                             // pio_Button:readdata -> pio_Button_s1_translator:av_readdata
	wire   [7:0] lcd_control_slave_translator_avalon_anti_slave_0_writedata;                                        // lcd_control_slave_translator:av_writedata -> lcd:writedata
	wire   [1:0] lcd_control_slave_translator_avalon_anti_slave_0_address;                                          // lcd_control_slave_translator:av_address -> lcd:address
	wire         lcd_control_slave_translator_avalon_anti_slave_0_write;                                            // lcd_control_slave_translator:av_write -> lcd:write
	wire         lcd_control_slave_translator_avalon_anti_slave_0_read;                                             // lcd_control_slave_translator:av_read -> lcd:read
	wire   [7:0] lcd_control_slave_translator_avalon_anti_slave_0_readdata;                                         // lcd:readdata -> lcd_control_slave_translator:av_readdata
	wire         lcd_control_slave_translator_avalon_anti_slave_0_begintransfer;                                    // lcd_control_slave_translator:av_begintransfer -> lcd:begintransfer
	wire  [15:0] uart_s1_translator_avalon_anti_slave_0_writedata;                                                  // uart_s1_translator:av_writedata -> uart:writedata
	wire   [2:0] uart_s1_translator_avalon_anti_slave_0_address;                                                    // uart_s1_translator:av_address -> uart:address
	wire         uart_s1_translator_avalon_anti_slave_0_chipselect;                                                 // uart_s1_translator:av_chipselect -> uart:chipselect
	wire         uart_s1_translator_avalon_anti_slave_0_write;                                                      // uart_s1_translator:av_write -> uart:write_n
	wire         uart_s1_translator_avalon_anti_slave_0_read;                                                       // uart_s1_translator:av_read -> uart:read_n
	wire  [15:0] uart_s1_translator_avalon_anti_slave_0_readdata;                                                   // uart:readdata -> uart_s1_translator:av_readdata
	wire         uart_s1_translator_avalon_anti_slave_0_begintransfer;                                              // uart_s1_translator:av_begintransfer -> uart:begintransfer
	wire  [15:0] timer_0_s1_translator_avalon_anti_slave_0_writedata;                                               // timer_0_s1_translator:av_writedata -> timer_0:writedata
	wire   [2:0] timer_0_s1_translator_avalon_anti_slave_0_address;                                                 // timer_0_s1_translator:av_address -> timer_0:address
	wire         timer_0_s1_translator_avalon_anti_slave_0_chipselect;                                              // timer_0_s1_translator:av_chipselect -> timer_0:chipselect
	wire         timer_0_s1_translator_avalon_anti_slave_0_write;                                                   // timer_0_s1_translator:av_write -> timer_0:write_n
	wire  [15:0] timer_0_s1_translator_avalon_anti_slave_0_readdata;                                                // timer_0:readdata -> timer_0_s1_translator:av_readdata
	wire   [1:0] pio_data_s1_translator_avalon_anti_slave_0_address;                                                // pio_Data_s1_translator:av_address -> pio_Data:address
	wire  [31:0] pio_data_s1_translator_avalon_anti_slave_0_readdata;                                               // pio_Data:readdata -> pio_Data_s1_translator:av_readdata
	wire  [31:0] pio_rdydata_s1_translator_avalon_anti_slave_0_writedata;                                           // pio_RdyData_s1_translator:av_writedata -> pio_RdyData:writedata
	wire   [1:0] pio_rdydata_s1_translator_avalon_anti_slave_0_address;                                             // pio_RdyData_s1_translator:av_address -> pio_RdyData:address
	wire         pio_rdydata_s1_translator_avalon_anti_slave_0_chipselect;                                          // pio_RdyData_s1_translator:av_chipselect -> pio_RdyData:chipselect
	wire         pio_rdydata_s1_translator_avalon_anti_slave_0_write;                                               // pio_RdyData_s1_translator:av_write -> pio_RdyData:write_n
	wire  [31:0] pio_rdydata_s1_translator_avalon_anti_slave_0_readdata;                                            // pio_RdyData:readdata -> pio_RdyData_s1_translator:av_readdata
	wire  [31:0] pio_dataread_s1_translator_avalon_anti_slave_0_writedata;                                          // pio_DataRead_s1_translator:av_writedata -> pio_DataRead:writedata
	wire   [2:0] pio_dataread_s1_translator_avalon_anti_slave_0_address;                                            // pio_DataRead_s1_translator:av_address -> pio_DataRead:address
	wire         pio_dataread_s1_translator_avalon_anti_slave_0_chipselect;                                         // pio_DataRead_s1_translator:av_chipselect -> pio_DataRead:chipselect
	wire         pio_dataread_s1_translator_avalon_anti_slave_0_write;                                              // pio_DataRead_s1_translator:av_write -> pio_DataRead:write_n
	wire  [31:0] pio_dataread_s1_translator_avalon_anti_slave_0_readdata;                                           // pio_DataRead:readdata -> pio_DataRead_s1_translator:av_readdata
	wire         uart_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest;                                  // uart_s1_translator:uav_waitrequest -> uart_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire   [2:0] uart_s1_translator_avalon_universal_slave_0_agent_m0_burstcount;                                   // uart_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> uart_s1_translator:uav_burstcount
	wire  [31:0] uart_s1_translator_avalon_universal_slave_0_agent_m0_writedata;                                    // uart_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> uart_s1_translator:uav_writedata
	wire  [18:0] uart_s1_translator_avalon_universal_slave_0_agent_m0_address;                                      // uart_s1_translator_avalon_universal_slave_0_agent:m0_address -> uart_s1_translator:uav_address
	wire         uart_s1_translator_avalon_universal_slave_0_agent_m0_write;                                        // uart_s1_translator_avalon_universal_slave_0_agent:m0_write -> uart_s1_translator:uav_write
	wire         uart_s1_translator_avalon_universal_slave_0_agent_m0_lock;                                         // uart_s1_translator_avalon_universal_slave_0_agent:m0_lock -> uart_s1_translator:uav_lock
	wire         uart_s1_translator_avalon_universal_slave_0_agent_m0_read;                                         // uart_s1_translator_avalon_universal_slave_0_agent:m0_read -> uart_s1_translator:uav_read
	wire  [31:0] uart_s1_translator_avalon_universal_slave_0_agent_m0_readdata;                                     // uart_s1_translator:uav_readdata -> uart_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	wire         uart_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                                // uart_s1_translator:uav_readdatavalid -> uart_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire         uart_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess;                                  // uart_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> uart_s1_translator:uav_debugaccess
	wire   [3:0] uart_s1_translator_avalon_universal_slave_0_agent_m0_byteenable;                                   // uart_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> uart_s1_translator:uav_byteenable
	wire         uart_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                           // uart_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> uart_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire         uart_s1_translator_avalon_universal_slave_0_agent_rf_source_valid;                                 // uart_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> uart_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire         uart_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                         // uart_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> uart_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [76:0] uart_s1_translator_avalon_universal_slave_0_agent_rf_source_data;                                  // uart_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> uart_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire         uart_s1_translator_avalon_universal_slave_0_agent_rf_source_ready;                                 // uart_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> uart_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire         uart_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                        // uart_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> uart_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire         uart_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                              // uart_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> uart_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire         uart_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;                      // uart_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> uart_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [76:0] uart_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                               // uart_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> uart_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire         uart_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                              // uart_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> uart_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire         uart_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                            // uart_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> uart_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire  [31:0] uart_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                             // uart_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> uart_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire         uart_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                            // uart_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> uart_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire         pio_dataread_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest;                          // pio_DataRead_s1_translator:uav_waitrequest -> pio_DataRead_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire   [2:0] pio_dataread_s1_translator_avalon_universal_slave_0_agent_m0_burstcount;                           // pio_DataRead_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> pio_DataRead_s1_translator:uav_burstcount
	wire  [31:0] pio_dataread_s1_translator_avalon_universal_slave_0_agent_m0_writedata;                            // pio_DataRead_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> pio_DataRead_s1_translator:uav_writedata
	wire  [18:0] pio_dataread_s1_translator_avalon_universal_slave_0_agent_m0_address;                              // pio_DataRead_s1_translator_avalon_universal_slave_0_agent:m0_address -> pio_DataRead_s1_translator:uav_address
	wire         pio_dataread_s1_translator_avalon_universal_slave_0_agent_m0_write;                                // pio_DataRead_s1_translator_avalon_universal_slave_0_agent:m0_write -> pio_DataRead_s1_translator:uav_write
	wire         pio_dataread_s1_translator_avalon_universal_slave_0_agent_m0_lock;                                 // pio_DataRead_s1_translator_avalon_universal_slave_0_agent:m0_lock -> pio_DataRead_s1_translator:uav_lock
	wire         pio_dataread_s1_translator_avalon_universal_slave_0_agent_m0_read;                                 // pio_DataRead_s1_translator_avalon_universal_slave_0_agent:m0_read -> pio_DataRead_s1_translator:uav_read
	wire  [31:0] pio_dataread_s1_translator_avalon_universal_slave_0_agent_m0_readdata;                             // pio_DataRead_s1_translator:uav_readdata -> pio_DataRead_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	wire         pio_dataread_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                        // pio_DataRead_s1_translator:uav_readdatavalid -> pio_DataRead_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire         pio_dataread_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess;                          // pio_DataRead_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> pio_DataRead_s1_translator:uav_debugaccess
	wire   [3:0] pio_dataread_s1_translator_avalon_universal_slave_0_agent_m0_byteenable;                           // pio_DataRead_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> pio_DataRead_s1_translator:uav_byteenable
	wire         pio_dataread_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                   // pio_DataRead_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> pio_DataRead_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire         pio_dataread_s1_translator_avalon_universal_slave_0_agent_rf_source_valid;                         // pio_DataRead_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> pio_DataRead_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire         pio_dataread_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                 // pio_DataRead_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> pio_DataRead_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [76:0] pio_dataread_s1_translator_avalon_universal_slave_0_agent_rf_source_data;                          // pio_DataRead_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> pio_DataRead_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire         pio_dataread_s1_translator_avalon_universal_slave_0_agent_rf_source_ready;                         // pio_DataRead_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> pio_DataRead_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire         pio_dataread_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                // pio_DataRead_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> pio_DataRead_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire         pio_dataread_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                      // pio_DataRead_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> pio_DataRead_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire         pio_dataread_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;              // pio_DataRead_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> pio_DataRead_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [76:0] pio_dataread_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                       // pio_DataRead_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> pio_DataRead_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire         pio_dataread_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                      // pio_DataRead_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> pio_DataRead_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire         pio_dataread_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                    // pio_DataRead_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> pio_DataRead_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire  [31:0] pio_dataread_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                     // pio_DataRead_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> pio_DataRead_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire         pio_dataread_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                    // pio_DataRead_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> pio_DataRead_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire         pio_rdydata_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest;                           // pio_RdyData_s1_translator:uav_waitrequest -> pio_RdyData_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire   [2:0] pio_rdydata_s1_translator_avalon_universal_slave_0_agent_m0_burstcount;                            // pio_RdyData_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> pio_RdyData_s1_translator:uav_burstcount
	wire  [31:0] pio_rdydata_s1_translator_avalon_universal_slave_0_agent_m0_writedata;                             // pio_RdyData_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> pio_RdyData_s1_translator:uav_writedata
	wire  [18:0] pio_rdydata_s1_translator_avalon_universal_slave_0_agent_m0_address;                               // pio_RdyData_s1_translator_avalon_universal_slave_0_agent:m0_address -> pio_RdyData_s1_translator:uav_address
	wire         pio_rdydata_s1_translator_avalon_universal_slave_0_agent_m0_write;                                 // pio_RdyData_s1_translator_avalon_universal_slave_0_agent:m0_write -> pio_RdyData_s1_translator:uav_write
	wire         pio_rdydata_s1_translator_avalon_universal_slave_0_agent_m0_lock;                                  // pio_RdyData_s1_translator_avalon_universal_slave_0_agent:m0_lock -> pio_RdyData_s1_translator:uav_lock
	wire         pio_rdydata_s1_translator_avalon_universal_slave_0_agent_m0_read;                                  // pio_RdyData_s1_translator_avalon_universal_slave_0_agent:m0_read -> pio_RdyData_s1_translator:uav_read
	wire  [31:0] pio_rdydata_s1_translator_avalon_universal_slave_0_agent_m0_readdata;                              // pio_RdyData_s1_translator:uav_readdata -> pio_RdyData_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	wire         pio_rdydata_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                         // pio_RdyData_s1_translator:uav_readdatavalid -> pio_RdyData_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire         pio_rdydata_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess;                           // pio_RdyData_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> pio_RdyData_s1_translator:uav_debugaccess
	wire   [3:0] pio_rdydata_s1_translator_avalon_universal_slave_0_agent_m0_byteenable;                            // pio_RdyData_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> pio_RdyData_s1_translator:uav_byteenable
	wire         pio_rdydata_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                    // pio_RdyData_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> pio_RdyData_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire         pio_rdydata_s1_translator_avalon_universal_slave_0_agent_rf_source_valid;                          // pio_RdyData_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> pio_RdyData_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire         pio_rdydata_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                  // pio_RdyData_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> pio_RdyData_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [76:0] pio_rdydata_s1_translator_avalon_universal_slave_0_agent_rf_source_data;                           // pio_RdyData_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> pio_RdyData_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire         pio_rdydata_s1_translator_avalon_universal_slave_0_agent_rf_source_ready;                          // pio_RdyData_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> pio_RdyData_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire         pio_rdydata_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                 // pio_RdyData_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> pio_RdyData_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire         pio_rdydata_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                       // pio_RdyData_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> pio_RdyData_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire         pio_rdydata_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;               // pio_RdyData_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> pio_RdyData_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [76:0] pio_rdydata_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                        // pio_RdyData_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> pio_RdyData_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire         pio_rdydata_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                       // pio_RdyData_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> pio_RdyData_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire         pio_rdydata_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                     // pio_RdyData_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> pio_RdyData_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire  [31:0] pio_rdydata_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                      // pio_RdyData_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> pio_RdyData_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire         pio_rdydata_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                     // pio_RdyData_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> pio_RdyData_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire         jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest;              // jtag_uart_avalon_jtag_slave_translator:uav_waitrequest -> jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire   [2:0] jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_burstcount;               // jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_burstcount -> jtag_uart_avalon_jtag_slave_translator:uav_burstcount
	wire  [31:0] jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_writedata;                // jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_writedata -> jtag_uart_avalon_jtag_slave_translator:uav_writedata
	wire  [18:0] jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_address;                  // jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_address -> jtag_uart_avalon_jtag_slave_translator:uav_address
	wire         jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_write;                    // jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_write -> jtag_uart_avalon_jtag_slave_translator:uav_write
	wire         jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_lock;                     // jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_lock -> jtag_uart_avalon_jtag_slave_translator:uav_lock
	wire         jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_read;                     // jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_read -> jtag_uart_avalon_jtag_slave_translator:uav_read
	wire  [31:0] jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_readdata;                 // jtag_uart_avalon_jtag_slave_translator:uav_readdata -> jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_readdata
	wire         jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid;            // jtag_uart_avalon_jtag_slave_translator:uav_readdatavalid -> jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire         jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess;              // jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_debugaccess -> jtag_uart_avalon_jtag_slave_translator:uav_debugaccess
	wire   [3:0] jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_byteenable;               // jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_byteenable -> jtag_uart_avalon_jtag_slave_translator:uav_byteenable
	wire         jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;       // jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire         jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_valid;             // jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_source_valid -> jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire         jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;     // jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [76:0] jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_data;              // jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_source_data -> jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire         jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_ready;             // jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire         jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;    // jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire         jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;          // jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire         jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;  // jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [76:0] jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;           // jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire         jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;          // jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_sink_ready -> jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire         jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;        // jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire  [31:0] jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;         // jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire         jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;        // jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire         lcd_control_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest;                        // lcd_control_slave_translator:uav_waitrequest -> lcd_control_slave_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire   [2:0] lcd_control_slave_translator_avalon_universal_slave_0_agent_m0_burstcount;                         // lcd_control_slave_translator_avalon_universal_slave_0_agent:m0_burstcount -> lcd_control_slave_translator:uav_burstcount
	wire  [31:0] lcd_control_slave_translator_avalon_universal_slave_0_agent_m0_writedata;                          // lcd_control_slave_translator_avalon_universal_slave_0_agent:m0_writedata -> lcd_control_slave_translator:uav_writedata
	wire  [18:0] lcd_control_slave_translator_avalon_universal_slave_0_agent_m0_address;                            // lcd_control_slave_translator_avalon_universal_slave_0_agent:m0_address -> lcd_control_slave_translator:uav_address
	wire         lcd_control_slave_translator_avalon_universal_slave_0_agent_m0_write;                              // lcd_control_slave_translator_avalon_universal_slave_0_agent:m0_write -> lcd_control_slave_translator:uav_write
	wire         lcd_control_slave_translator_avalon_universal_slave_0_agent_m0_lock;                               // lcd_control_slave_translator_avalon_universal_slave_0_agent:m0_lock -> lcd_control_slave_translator:uav_lock
	wire         lcd_control_slave_translator_avalon_universal_slave_0_agent_m0_read;                               // lcd_control_slave_translator_avalon_universal_slave_0_agent:m0_read -> lcd_control_slave_translator:uav_read
	wire  [31:0] lcd_control_slave_translator_avalon_universal_slave_0_agent_m0_readdata;                           // lcd_control_slave_translator:uav_readdata -> lcd_control_slave_translator_avalon_universal_slave_0_agent:m0_readdata
	wire         lcd_control_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                      // lcd_control_slave_translator:uav_readdatavalid -> lcd_control_slave_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire         lcd_control_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess;                        // lcd_control_slave_translator_avalon_universal_slave_0_agent:m0_debugaccess -> lcd_control_slave_translator:uav_debugaccess
	wire   [3:0] lcd_control_slave_translator_avalon_universal_slave_0_agent_m0_byteenable;                         // lcd_control_slave_translator_avalon_universal_slave_0_agent:m0_byteenable -> lcd_control_slave_translator:uav_byteenable
	wire         lcd_control_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                 // lcd_control_slave_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> lcd_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire         lcd_control_slave_translator_avalon_universal_slave_0_agent_rf_source_valid;                       // lcd_control_slave_translator_avalon_universal_slave_0_agent:rf_source_valid -> lcd_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire         lcd_control_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;               // lcd_control_slave_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> lcd_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [76:0] lcd_control_slave_translator_avalon_universal_slave_0_agent_rf_source_data;                        // lcd_control_slave_translator_avalon_universal_slave_0_agent:rf_source_data -> lcd_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire         lcd_control_slave_translator_avalon_universal_slave_0_agent_rf_source_ready;                       // lcd_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> lcd_control_slave_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire         lcd_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;              // lcd_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> lcd_control_slave_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire         lcd_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                    // lcd_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> lcd_control_slave_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire         lcd_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;            // lcd_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> lcd_control_slave_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [76:0] lcd_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                     // lcd_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> lcd_control_slave_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire         lcd_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                    // lcd_control_slave_translator_avalon_universal_slave_0_agent:rf_sink_ready -> lcd_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire         lcd_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                  // lcd_control_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> lcd_control_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire  [31:0] lcd_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                   // lcd_control_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> lcd_control_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire         lcd_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                  // lcd_control_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> lcd_control_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire         pio_ledr_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest;                              // pio_LEDR_s1_translator:uav_waitrequest -> pio_LEDR_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire   [2:0] pio_ledr_s1_translator_avalon_universal_slave_0_agent_m0_burstcount;                               // pio_LEDR_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> pio_LEDR_s1_translator:uav_burstcount
	wire  [31:0] pio_ledr_s1_translator_avalon_universal_slave_0_agent_m0_writedata;                                // pio_LEDR_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> pio_LEDR_s1_translator:uav_writedata
	wire  [18:0] pio_ledr_s1_translator_avalon_universal_slave_0_agent_m0_address;                                  // pio_LEDR_s1_translator_avalon_universal_slave_0_agent:m0_address -> pio_LEDR_s1_translator:uav_address
	wire         pio_ledr_s1_translator_avalon_universal_slave_0_agent_m0_write;                                    // pio_LEDR_s1_translator_avalon_universal_slave_0_agent:m0_write -> pio_LEDR_s1_translator:uav_write
	wire         pio_ledr_s1_translator_avalon_universal_slave_0_agent_m0_lock;                                     // pio_LEDR_s1_translator_avalon_universal_slave_0_agent:m0_lock -> pio_LEDR_s1_translator:uav_lock
	wire         pio_ledr_s1_translator_avalon_universal_slave_0_agent_m0_read;                                     // pio_LEDR_s1_translator_avalon_universal_slave_0_agent:m0_read -> pio_LEDR_s1_translator:uav_read
	wire  [31:0] pio_ledr_s1_translator_avalon_universal_slave_0_agent_m0_readdata;                                 // pio_LEDR_s1_translator:uav_readdata -> pio_LEDR_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	wire         pio_ledr_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                            // pio_LEDR_s1_translator:uav_readdatavalid -> pio_LEDR_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire         pio_ledr_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess;                              // pio_LEDR_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> pio_LEDR_s1_translator:uav_debugaccess
	wire   [3:0] pio_ledr_s1_translator_avalon_universal_slave_0_agent_m0_byteenable;                               // pio_LEDR_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> pio_LEDR_s1_translator:uav_byteenable
	wire         pio_ledr_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                       // pio_LEDR_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> pio_LEDR_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire         pio_ledr_s1_translator_avalon_universal_slave_0_agent_rf_source_valid;                             // pio_LEDR_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> pio_LEDR_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire         pio_ledr_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                     // pio_LEDR_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> pio_LEDR_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [76:0] pio_ledr_s1_translator_avalon_universal_slave_0_agent_rf_source_data;                              // pio_LEDR_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> pio_LEDR_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire         pio_ledr_s1_translator_avalon_universal_slave_0_agent_rf_source_ready;                             // pio_LEDR_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> pio_LEDR_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire         pio_ledr_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                    // pio_LEDR_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> pio_LEDR_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire         pio_ledr_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                          // pio_LEDR_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> pio_LEDR_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire         pio_ledr_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;                  // pio_LEDR_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> pio_LEDR_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [76:0] pio_ledr_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                           // pio_LEDR_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> pio_LEDR_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire         pio_ledr_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                          // pio_LEDR_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> pio_LEDR_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire         pio_ledr_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                        // pio_LEDR_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> pio_LEDR_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire  [31:0] pio_ledr_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                         // pio_LEDR_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> pio_LEDR_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire         pio_ledr_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                        // pio_LEDR_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> pio_LEDR_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire         nios2_qsys_instruction_master_translator_avalon_universal_master_0_waitrequest;                    // nios2_qsys_instruction_master_translator_avalon_universal_master_0_agent:av_waitrequest -> nios2_qsys_instruction_master_translator:uav_waitrequest
	wire   [2:0] nios2_qsys_instruction_master_translator_avalon_universal_master_0_burstcount;                     // nios2_qsys_instruction_master_translator:uav_burstcount -> nios2_qsys_instruction_master_translator_avalon_universal_master_0_agent:av_burstcount
	wire  [31:0] nios2_qsys_instruction_master_translator_avalon_universal_master_0_writedata;                      // nios2_qsys_instruction_master_translator:uav_writedata -> nios2_qsys_instruction_master_translator_avalon_universal_master_0_agent:av_writedata
	wire  [18:0] nios2_qsys_instruction_master_translator_avalon_universal_master_0_address;                        // nios2_qsys_instruction_master_translator:uav_address -> nios2_qsys_instruction_master_translator_avalon_universal_master_0_agent:av_address
	wire         nios2_qsys_instruction_master_translator_avalon_universal_master_0_lock;                           // nios2_qsys_instruction_master_translator:uav_lock -> nios2_qsys_instruction_master_translator_avalon_universal_master_0_agent:av_lock
	wire         nios2_qsys_instruction_master_translator_avalon_universal_master_0_write;                          // nios2_qsys_instruction_master_translator:uav_write -> nios2_qsys_instruction_master_translator_avalon_universal_master_0_agent:av_write
	wire         nios2_qsys_instruction_master_translator_avalon_universal_master_0_read;                           // nios2_qsys_instruction_master_translator:uav_read -> nios2_qsys_instruction_master_translator_avalon_universal_master_0_agent:av_read
	wire  [31:0] nios2_qsys_instruction_master_translator_avalon_universal_master_0_readdata;                       // nios2_qsys_instruction_master_translator_avalon_universal_master_0_agent:av_readdata -> nios2_qsys_instruction_master_translator:uav_readdata
	wire         nios2_qsys_instruction_master_translator_avalon_universal_master_0_debugaccess;                    // nios2_qsys_instruction_master_translator:uav_debugaccess -> nios2_qsys_instruction_master_translator_avalon_universal_master_0_agent:av_debugaccess
	wire   [3:0] nios2_qsys_instruction_master_translator_avalon_universal_master_0_byteenable;                     // nios2_qsys_instruction_master_translator:uav_byteenable -> nios2_qsys_instruction_master_translator_avalon_universal_master_0_agent:av_byteenable
	wire         nios2_qsys_instruction_master_translator_avalon_universal_master_0_readdatavalid;                  // nios2_qsys_instruction_master_translator_avalon_universal_master_0_agent:av_readdatavalid -> nios2_qsys_instruction_master_translator:uav_readdatavalid
	wire         nios2_qsys_data_master_translator_avalon_universal_master_0_waitrequest;                           // nios2_qsys_data_master_translator_avalon_universal_master_0_agent:av_waitrequest -> nios2_qsys_data_master_translator:uav_waitrequest
	wire   [2:0] nios2_qsys_data_master_translator_avalon_universal_master_0_burstcount;                            // nios2_qsys_data_master_translator:uav_burstcount -> nios2_qsys_data_master_translator_avalon_universal_master_0_agent:av_burstcount
	wire  [31:0] nios2_qsys_data_master_translator_avalon_universal_master_0_writedata;                             // nios2_qsys_data_master_translator:uav_writedata -> nios2_qsys_data_master_translator_avalon_universal_master_0_agent:av_writedata
	wire  [18:0] nios2_qsys_data_master_translator_avalon_universal_master_0_address;                               // nios2_qsys_data_master_translator:uav_address -> nios2_qsys_data_master_translator_avalon_universal_master_0_agent:av_address
	wire         nios2_qsys_data_master_translator_avalon_universal_master_0_lock;                                  // nios2_qsys_data_master_translator:uav_lock -> nios2_qsys_data_master_translator_avalon_universal_master_0_agent:av_lock
	wire         nios2_qsys_data_master_translator_avalon_universal_master_0_write;                                 // nios2_qsys_data_master_translator:uav_write -> nios2_qsys_data_master_translator_avalon_universal_master_0_agent:av_write
	wire         nios2_qsys_data_master_translator_avalon_universal_master_0_read;                                  // nios2_qsys_data_master_translator:uav_read -> nios2_qsys_data_master_translator_avalon_universal_master_0_agent:av_read
	wire  [31:0] nios2_qsys_data_master_translator_avalon_universal_master_0_readdata;                              // nios2_qsys_data_master_translator_avalon_universal_master_0_agent:av_readdata -> nios2_qsys_data_master_translator:uav_readdata
	wire         nios2_qsys_data_master_translator_avalon_universal_master_0_debugaccess;                           // nios2_qsys_data_master_translator:uav_debugaccess -> nios2_qsys_data_master_translator_avalon_universal_master_0_agent:av_debugaccess
	wire   [3:0] nios2_qsys_data_master_translator_avalon_universal_master_0_byteenable;                            // nios2_qsys_data_master_translator:uav_byteenable -> nios2_qsys_data_master_translator_avalon_universal_master_0_agent:av_byteenable
	wire         nios2_qsys_data_master_translator_avalon_universal_master_0_readdatavalid;                         // nios2_qsys_data_master_translator_avalon_universal_master_0_agent:av_readdatavalid -> nios2_qsys_data_master_translator:uav_readdatavalid
	wire         onchip_memory_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest;                         // onchip_memory_s1_translator:uav_waitrequest -> onchip_memory_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire   [2:0] onchip_memory_s1_translator_avalon_universal_slave_0_agent_m0_burstcount;                          // onchip_memory_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> onchip_memory_s1_translator:uav_burstcount
	wire  [31:0] onchip_memory_s1_translator_avalon_universal_slave_0_agent_m0_writedata;                           // onchip_memory_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> onchip_memory_s1_translator:uav_writedata
	wire  [18:0] onchip_memory_s1_translator_avalon_universal_slave_0_agent_m0_address;                             // onchip_memory_s1_translator_avalon_universal_slave_0_agent:m0_address -> onchip_memory_s1_translator:uav_address
	wire         onchip_memory_s1_translator_avalon_universal_slave_0_agent_m0_write;                               // onchip_memory_s1_translator_avalon_universal_slave_0_agent:m0_write -> onchip_memory_s1_translator:uav_write
	wire         onchip_memory_s1_translator_avalon_universal_slave_0_agent_m0_lock;                                // onchip_memory_s1_translator_avalon_universal_slave_0_agent:m0_lock -> onchip_memory_s1_translator:uav_lock
	wire         onchip_memory_s1_translator_avalon_universal_slave_0_agent_m0_read;                                // onchip_memory_s1_translator_avalon_universal_slave_0_agent:m0_read -> onchip_memory_s1_translator:uav_read
	wire  [31:0] onchip_memory_s1_translator_avalon_universal_slave_0_agent_m0_readdata;                            // onchip_memory_s1_translator:uav_readdata -> onchip_memory_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	wire         onchip_memory_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                       // onchip_memory_s1_translator:uav_readdatavalid -> onchip_memory_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire         onchip_memory_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess;                         // onchip_memory_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> onchip_memory_s1_translator:uav_debugaccess
	wire   [3:0] onchip_memory_s1_translator_avalon_universal_slave_0_agent_m0_byteenable;                          // onchip_memory_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> onchip_memory_s1_translator:uav_byteenable
	wire         onchip_memory_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                  // onchip_memory_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> onchip_memory_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire         onchip_memory_s1_translator_avalon_universal_slave_0_agent_rf_source_valid;                        // onchip_memory_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> onchip_memory_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire         onchip_memory_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                // onchip_memory_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> onchip_memory_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [76:0] onchip_memory_s1_translator_avalon_universal_slave_0_agent_rf_source_data;                         // onchip_memory_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> onchip_memory_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire         onchip_memory_s1_translator_avalon_universal_slave_0_agent_rf_source_ready;                        // onchip_memory_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> onchip_memory_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire         onchip_memory_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;               // onchip_memory_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> onchip_memory_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire         onchip_memory_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                     // onchip_memory_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> onchip_memory_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire         onchip_memory_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;             // onchip_memory_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> onchip_memory_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [76:0] onchip_memory_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                      // onchip_memory_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> onchip_memory_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire         onchip_memory_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                     // onchip_memory_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> onchip_memory_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire         onchip_memory_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                   // onchip_memory_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> onchip_memory_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire  [31:0] onchip_memory_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                    // onchip_memory_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> onchip_memory_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire         onchip_memory_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                   // onchip_memory_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> onchip_memory_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire         pio_sw_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest;                                // pio_SW_s1_translator:uav_waitrequest -> pio_SW_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire   [2:0] pio_sw_s1_translator_avalon_universal_slave_0_agent_m0_burstcount;                                 // pio_SW_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> pio_SW_s1_translator:uav_burstcount
	wire  [31:0] pio_sw_s1_translator_avalon_universal_slave_0_agent_m0_writedata;                                  // pio_SW_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> pio_SW_s1_translator:uav_writedata
	wire  [18:0] pio_sw_s1_translator_avalon_universal_slave_0_agent_m0_address;                                    // pio_SW_s1_translator_avalon_universal_slave_0_agent:m0_address -> pio_SW_s1_translator:uav_address
	wire         pio_sw_s1_translator_avalon_universal_slave_0_agent_m0_write;                                      // pio_SW_s1_translator_avalon_universal_slave_0_agent:m0_write -> pio_SW_s1_translator:uav_write
	wire         pio_sw_s1_translator_avalon_universal_slave_0_agent_m0_lock;                                       // pio_SW_s1_translator_avalon_universal_slave_0_agent:m0_lock -> pio_SW_s1_translator:uav_lock
	wire         pio_sw_s1_translator_avalon_universal_slave_0_agent_m0_read;                                       // pio_SW_s1_translator_avalon_universal_slave_0_agent:m0_read -> pio_SW_s1_translator:uav_read
	wire  [31:0] pio_sw_s1_translator_avalon_universal_slave_0_agent_m0_readdata;                                   // pio_SW_s1_translator:uav_readdata -> pio_SW_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	wire         pio_sw_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                              // pio_SW_s1_translator:uav_readdatavalid -> pio_SW_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire         pio_sw_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess;                                // pio_SW_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> pio_SW_s1_translator:uav_debugaccess
	wire   [3:0] pio_sw_s1_translator_avalon_universal_slave_0_agent_m0_byteenable;                                 // pio_SW_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> pio_SW_s1_translator:uav_byteenable
	wire         pio_sw_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                         // pio_SW_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> pio_SW_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire         pio_sw_s1_translator_avalon_universal_slave_0_agent_rf_source_valid;                               // pio_SW_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> pio_SW_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire         pio_sw_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                       // pio_SW_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> pio_SW_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [76:0] pio_sw_s1_translator_avalon_universal_slave_0_agent_rf_source_data;                                // pio_SW_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> pio_SW_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire         pio_sw_s1_translator_avalon_universal_slave_0_agent_rf_source_ready;                               // pio_SW_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> pio_SW_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire         pio_sw_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                      // pio_SW_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> pio_SW_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire         pio_sw_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                            // pio_SW_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> pio_SW_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire         pio_sw_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;                    // pio_SW_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> pio_SW_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [76:0] pio_sw_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                             // pio_SW_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> pio_SW_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire         pio_sw_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                            // pio_SW_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> pio_SW_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire         pio_sw_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                          // pio_SW_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> pio_SW_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire  [31:0] pio_sw_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                           // pio_SW_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> pio_SW_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire         pio_sw_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                          // pio_SW_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> pio_SW_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire         sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest;                 // sysid_qsys_control_slave_translator:uav_waitrequest -> sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire   [2:0] sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent_m0_burstcount;                  // sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent:m0_burstcount -> sysid_qsys_control_slave_translator:uav_burstcount
	wire  [31:0] sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent_m0_writedata;                   // sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent:m0_writedata -> sysid_qsys_control_slave_translator:uav_writedata
	wire  [18:0] sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent_m0_address;                     // sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent:m0_address -> sysid_qsys_control_slave_translator:uav_address
	wire         sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent_m0_write;                       // sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent:m0_write -> sysid_qsys_control_slave_translator:uav_write
	wire         sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent_m0_lock;                        // sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent:m0_lock -> sysid_qsys_control_slave_translator:uav_lock
	wire         sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent_m0_read;                        // sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent:m0_read -> sysid_qsys_control_slave_translator:uav_read
	wire  [31:0] sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent_m0_readdata;                    // sysid_qsys_control_slave_translator:uav_readdata -> sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent:m0_readdata
	wire         sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid;               // sysid_qsys_control_slave_translator:uav_readdatavalid -> sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire         sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess;                 // sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent:m0_debugaccess -> sysid_qsys_control_slave_translator:uav_debugaccess
	wire   [3:0] sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent_m0_byteenable;                  // sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent:m0_byteenable -> sysid_qsys_control_slave_translator:uav_byteenable
	wire         sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;          // sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire         sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent_rf_source_valid;                // sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent:rf_source_valid -> sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire         sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;        // sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [76:0] sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent_rf_source_data;                 // sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent:rf_source_data -> sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire         sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent_rf_source_ready;                // sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire         sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;       // sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire         sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;             // sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire         sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;     // sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [76:0] sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;              // sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire         sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;             // sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent:rf_sink_ready -> sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire         sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;           // sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire  [31:0] sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;            // sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire         sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;           // sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire         nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_waitrequest;             // nios2_qsys_jtag_debug_module_translator:uav_waitrequest -> nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire   [2:0] nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_burstcount;              // nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_burstcount -> nios2_qsys_jtag_debug_module_translator:uav_burstcount
	wire  [31:0] nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_writedata;               // nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_writedata -> nios2_qsys_jtag_debug_module_translator:uav_writedata
	wire  [18:0] nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_address;                 // nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_address -> nios2_qsys_jtag_debug_module_translator:uav_address
	wire         nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_write;                   // nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_write -> nios2_qsys_jtag_debug_module_translator:uav_write
	wire         nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_lock;                    // nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_lock -> nios2_qsys_jtag_debug_module_translator:uav_lock
	wire         nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_read;                    // nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_read -> nios2_qsys_jtag_debug_module_translator:uav_read
	wire  [31:0] nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_readdata;                // nios2_qsys_jtag_debug_module_translator:uav_readdata -> nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_readdata
	wire         nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_readdatavalid;           // nios2_qsys_jtag_debug_module_translator:uav_readdatavalid -> nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire         nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_debugaccess;             // nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_debugaccess -> nios2_qsys_jtag_debug_module_translator:uav_debugaccess
	wire   [3:0] nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_byteenable;              // nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_byteenable -> nios2_qsys_jtag_debug_module_translator:uav_byteenable
	wire         nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;      // nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire         nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_valid;            // nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_source_valid -> nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire         nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;    // nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [76:0] nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_data;             // nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_source_data -> nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire         nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_ready;            // nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire         nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;   // nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire         nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;         // nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire         nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket; // nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [76:0] nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;          // nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire         nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;         // nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_sink_ready -> nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire         nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;       // nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire  [31:0] nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;        // nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire         nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;       // nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire         pio_ledg_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest;                              // pio_LEDG_s1_translator:uav_waitrequest -> pio_LEDG_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire   [2:0] pio_ledg_s1_translator_avalon_universal_slave_0_agent_m0_burstcount;                               // pio_LEDG_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> pio_LEDG_s1_translator:uav_burstcount
	wire  [31:0] pio_ledg_s1_translator_avalon_universal_slave_0_agent_m0_writedata;                                // pio_LEDG_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> pio_LEDG_s1_translator:uav_writedata
	wire  [18:0] pio_ledg_s1_translator_avalon_universal_slave_0_agent_m0_address;                                  // pio_LEDG_s1_translator_avalon_universal_slave_0_agent:m0_address -> pio_LEDG_s1_translator:uav_address
	wire         pio_ledg_s1_translator_avalon_universal_slave_0_agent_m0_write;                                    // pio_LEDG_s1_translator_avalon_universal_slave_0_agent:m0_write -> pio_LEDG_s1_translator:uav_write
	wire         pio_ledg_s1_translator_avalon_universal_slave_0_agent_m0_lock;                                     // pio_LEDG_s1_translator_avalon_universal_slave_0_agent:m0_lock -> pio_LEDG_s1_translator:uav_lock
	wire         pio_ledg_s1_translator_avalon_universal_slave_0_agent_m0_read;                                     // pio_LEDG_s1_translator_avalon_universal_slave_0_agent:m0_read -> pio_LEDG_s1_translator:uav_read
	wire  [31:0] pio_ledg_s1_translator_avalon_universal_slave_0_agent_m0_readdata;                                 // pio_LEDG_s1_translator:uav_readdata -> pio_LEDG_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	wire         pio_ledg_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                            // pio_LEDG_s1_translator:uav_readdatavalid -> pio_LEDG_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire         pio_ledg_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess;                              // pio_LEDG_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> pio_LEDG_s1_translator:uav_debugaccess
	wire   [3:0] pio_ledg_s1_translator_avalon_universal_slave_0_agent_m0_byteenable;                               // pio_LEDG_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> pio_LEDG_s1_translator:uav_byteenable
	wire         pio_ledg_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                       // pio_LEDG_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> pio_LEDG_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire         pio_ledg_s1_translator_avalon_universal_slave_0_agent_rf_source_valid;                             // pio_LEDG_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> pio_LEDG_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire         pio_ledg_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                     // pio_LEDG_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> pio_LEDG_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [76:0] pio_ledg_s1_translator_avalon_universal_slave_0_agent_rf_source_data;                              // pio_LEDG_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> pio_LEDG_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire         pio_ledg_s1_translator_avalon_universal_slave_0_agent_rf_source_ready;                             // pio_LEDG_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> pio_LEDG_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire         pio_ledg_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                    // pio_LEDG_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> pio_LEDG_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire         pio_ledg_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                          // pio_LEDG_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> pio_LEDG_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire         pio_ledg_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;                  // pio_LEDG_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> pio_LEDG_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [76:0] pio_ledg_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                           // pio_LEDG_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> pio_LEDG_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire         pio_ledg_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                          // pio_LEDG_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> pio_LEDG_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire         pio_ledg_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                        // pio_LEDG_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> pio_LEDG_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire  [31:0] pio_ledg_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                         // pio_LEDG_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> pio_LEDG_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire         pio_ledg_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                        // pio_LEDG_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> pio_LEDG_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire         pio_data_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest;                              // pio_Data_s1_translator:uav_waitrequest -> pio_Data_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire   [2:0] pio_data_s1_translator_avalon_universal_slave_0_agent_m0_burstcount;                               // pio_Data_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> pio_Data_s1_translator:uav_burstcount
	wire  [31:0] pio_data_s1_translator_avalon_universal_slave_0_agent_m0_writedata;                                // pio_Data_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> pio_Data_s1_translator:uav_writedata
	wire  [18:0] pio_data_s1_translator_avalon_universal_slave_0_agent_m0_address;                                  // pio_Data_s1_translator_avalon_universal_slave_0_agent:m0_address -> pio_Data_s1_translator:uav_address
	wire         pio_data_s1_translator_avalon_universal_slave_0_agent_m0_write;                                    // pio_Data_s1_translator_avalon_universal_slave_0_agent:m0_write -> pio_Data_s1_translator:uav_write
	wire         pio_data_s1_translator_avalon_universal_slave_0_agent_m0_lock;                                     // pio_Data_s1_translator_avalon_universal_slave_0_agent:m0_lock -> pio_Data_s1_translator:uav_lock
	wire         pio_data_s1_translator_avalon_universal_slave_0_agent_m0_read;                                     // pio_Data_s1_translator_avalon_universal_slave_0_agent:m0_read -> pio_Data_s1_translator:uav_read
	wire  [31:0] pio_data_s1_translator_avalon_universal_slave_0_agent_m0_readdata;                                 // pio_Data_s1_translator:uav_readdata -> pio_Data_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	wire         pio_data_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                            // pio_Data_s1_translator:uav_readdatavalid -> pio_Data_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire         pio_data_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess;                              // pio_Data_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> pio_Data_s1_translator:uav_debugaccess
	wire   [3:0] pio_data_s1_translator_avalon_universal_slave_0_agent_m0_byteenable;                               // pio_Data_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> pio_Data_s1_translator:uav_byteenable
	wire         pio_data_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                       // pio_Data_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> pio_Data_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire         pio_data_s1_translator_avalon_universal_slave_0_agent_rf_source_valid;                             // pio_Data_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> pio_Data_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire         pio_data_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                     // pio_Data_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> pio_Data_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [76:0] pio_data_s1_translator_avalon_universal_slave_0_agent_rf_source_data;                              // pio_Data_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> pio_Data_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire         pio_data_s1_translator_avalon_universal_slave_0_agent_rf_source_ready;                             // pio_Data_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> pio_Data_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire         pio_data_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                    // pio_Data_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> pio_Data_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire         pio_data_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                          // pio_Data_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> pio_Data_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire         pio_data_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;                  // pio_Data_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> pio_Data_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [76:0] pio_data_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                           // pio_Data_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> pio_Data_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire         pio_data_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                          // pio_Data_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> pio_Data_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire         pio_data_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                        // pio_Data_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> pio_Data_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire  [31:0] pio_data_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                         // pio_Data_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> pio_Data_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire         pio_data_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                        // pio_Data_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> pio_Data_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire         pio_button_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest;                            // pio_Button_s1_translator:uav_waitrequest -> pio_Button_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire   [2:0] pio_button_s1_translator_avalon_universal_slave_0_agent_m0_burstcount;                             // pio_Button_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> pio_Button_s1_translator:uav_burstcount
	wire  [31:0] pio_button_s1_translator_avalon_universal_slave_0_agent_m0_writedata;                              // pio_Button_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> pio_Button_s1_translator:uav_writedata
	wire  [18:0] pio_button_s1_translator_avalon_universal_slave_0_agent_m0_address;                                // pio_Button_s1_translator_avalon_universal_slave_0_agent:m0_address -> pio_Button_s1_translator:uav_address
	wire         pio_button_s1_translator_avalon_universal_slave_0_agent_m0_write;                                  // pio_Button_s1_translator_avalon_universal_slave_0_agent:m0_write -> pio_Button_s1_translator:uav_write
	wire         pio_button_s1_translator_avalon_universal_slave_0_agent_m0_lock;                                   // pio_Button_s1_translator_avalon_universal_slave_0_agent:m0_lock -> pio_Button_s1_translator:uav_lock
	wire         pio_button_s1_translator_avalon_universal_slave_0_agent_m0_read;                                   // pio_Button_s1_translator_avalon_universal_slave_0_agent:m0_read -> pio_Button_s1_translator:uav_read
	wire  [31:0] pio_button_s1_translator_avalon_universal_slave_0_agent_m0_readdata;                               // pio_Button_s1_translator:uav_readdata -> pio_Button_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	wire         pio_button_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                          // pio_Button_s1_translator:uav_readdatavalid -> pio_Button_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire         pio_button_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess;                            // pio_Button_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> pio_Button_s1_translator:uav_debugaccess
	wire   [3:0] pio_button_s1_translator_avalon_universal_slave_0_agent_m0_byteenable;                             // pio_Button_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> pio_Button_s1_translator:uav_byteenable
	wire         pio_button_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                     // pio_Button_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> pio_Button_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire         pio_button_s1_translator_avalon_universal_slave_0_agent_rf_source_valid;                           // pio_Button_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> pio_Button_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire         pio_button_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                   // pio_Button_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> pio_Button_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [76:0] pio_button_s1_translator_avalon_universal_slave_0_agent_rf_source_data;                            // pio_Button_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> pio_Button_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire         pio_button_s1_translator_avalon_universal_slave_0_agent_rf_source_ready;                           // pio_Button_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> pio_Button_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire         pio_button_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                  // pio_Button_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> pio_Button_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire         pio_button_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                        // pio_Button_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> pio_Button_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire         pio_button_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;                // pio_Button_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> pio_Button_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [76:0] pio_button_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                         // pio_Button_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> pio_Button_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire         pio_button_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                        // pio_Button_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> pio_Button_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire         pio_button_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                      // pio_Button_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> pio_Button_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire  [31:0] pio_button_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                       // pio_Button_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> pio_Button_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire         pio_button_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                      // pio_Button_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> pio_Button_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire         timer_0_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest;                               // timer_0_s1_translator:uav_waitrequest -> timer_0_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire   [2:0] timer_0_s1_translator_avalon_universal_slave_0_agent_m0_burstcount;                                // timer_0_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> timer_0_s1_translator:uav_burstcount
	wire  [31:0] timer_0_s1_translator_avalon_universal_slave_0_agent_m0_writedata;                                 // timer_0_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> timer_0_s1_translator:uav_writedata
	wire  [18:0] timer_0_s1_translator_avalon_universal_slave_0_agent_m0_address;                                   // timer_0_s1_translator_avalon_universal_slave_0_agent:m0_address -> timer_0_s1_translator:uav_address
	wire         timer_0_s1_translator_avalon_universal_slave_0_agent_m0_write;                                     // timer_0_s1_translator_avalon_universal_slave_0_agent:m0_write -> timer_0_s1_translator:uav_write
	wire         timer_0_s1_translator_avalon_universal_slave_0_agent_m0_lock;                                      // timer_0_s1_translator_avalon_universal_slave_0_agent:m0_lock -> timer_0_s1_translator:uav_lock
	wire         timer_0_s1_translator_avalon_universal_slave_0_agent_m0_read;                                      // timer_0_s1_translator_avalon_universal_slave_0_agent:m0_read -> timer_0_s1_translator:uav_read
	wire  [31:0] timer_0_s1_translator_avalon_universal_slave_0_agent_m0_readdata;                                  // timer_0_s1_translator:uav_readdata -> timer_0_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	wire         timer_0_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                             // timer_0_s1_translator:uav_readdatavalid -> timer_0_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire         timer_0_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess;                               // timer_0_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> timer_0_s1_translator:uav_debugaccess
	wire   [3:0] timer_0_s1_translator_avalon_universal_slave_0_agent_m0_byteenable;                                // timer_0_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> timer_0_s1_translator:uav_byteenable
	wire         timer_0_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                        // timer_0_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> timer_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire         timer_0_s1_translator_avalon_universal_slave_0_agent_rf_source_valid;                              // timer_0_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> timer_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire         timer_0_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                      // timer_0_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> timer_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [76:0] timer_0_s1_translator_avalon_universal_slave_0_agent_rf_source_data;                               // timer_0_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> timer_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire         timer_0_s1_translator_avalon_universal_slave_0_agent_rf_source_ready;                              // timer_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> timer_0_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire         timer_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                     // timer_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> timer_0_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire         timer_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                           // timer_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> timer_0_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire         timer_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;                   // timer_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> timer_0_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [76:0] timer_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                            // timer_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> timer_0_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire         timer_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                           // timer_0_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> timer_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire         timer_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                         // timer_0_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> timer_0_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire  [31:0] timer_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                          // timer_0_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> timer_0_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire         timer_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                         // timer_0_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> timer_0_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire         nios2_qsys_instruction_master_translator_avalon_universal_master_0_agent_cp_endofpacket;           // nios2_qsys_instruction_master_translator_avalon_universal_master_0_agent:cp_endofpacket -> addr_router:sink_endofpacket
	wire         nios2_qsys_instruction_master_translator_avalon_universal_master_0_agent_cp_valid;                 // nios2_qsys_instruction_master_translator_avalon_universal_master_0_agent:cp_valid -> addr_router:sink_valid
	wire         nios2_qsys_instruction_master_translator_avalon_universal_master_0_agent_cp_startofpacket;         // nios2_qsys_instruction_master_translator_avalon_universal_master_0_agent:cp_startofpacket -> addr_router:sink_startofpacket
	wire  [75:0] nios2_qsys_instruction_master_translator_avalon_universal_master_0_agent_cp_data;                  // nios2_qsys_instruction_master_translator_avalon_universal_master_0_agent:cp_data -> addr_router:sink_data
	wire         nios2_qsys_instruction_master_translator_avalon_universal_master_0_agent_cp_ready;                 // addr_router:sink_ready -> nios2_qsys_instruction_master_translator_avalon_universal_master_0_agent:cp_ready
	wire         nios2_qsys_data_master_translator_avalon_universal_master_0_agent_cp_endofpacket;                  // nios2_qsys_data_master_translator_avalon_universal_master_0_agent:cp_endofpacket -> addr_router_001:sink_endofpacket
	wire         nios2_qsys_data_master_translator_avalon_universal_master_0_agent_cp_valid;                        // nios2_qsys_data_master_translator_avalon_universal_master_0_agent:cp_valid -> addr_router_001:sink_valid
	wire         nios2_qsys_data_master_translator_avalon_universal_master_0_agent_cp_startofpacket;                // nios2_qsys_data_master_translator_avalon_universal_master_0_agent:cp_startofpacket -> addr_router_001:sink_startofpacket
	wire  [75:0] nios2_qsys_data_master_translator_avalon_universal_master_0_agent_cp_data;                         // nios2_qsys_data_master_translator_avalon_universal_master_0_agent:cp_data -> addr_router_001:sink_data
	wire         nios2_qsys_data_master_translator_avalon_universal_master_0_agent_cp_ready;                        // addr_router_001:sink_ready -> nios2_qsys_data_master_translator_avalon_universal_master_0_agent:cp_ready
	wire         nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_endofpacket;             // nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router:sink_endofpacket
	wire         nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_valid;                   // nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent:rp_valid -> id_router:sink_valid
	wire         nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_startofpacket;           // nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router:sink_startofpacket
	wire  [75:0] nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_data;                    // nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent:rp_data -> id_router:sink_data
	wire         nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_ready;                   // id_router:sink_ready -> nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent:rp_ready
	wire         onchip_memory_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket;                         // onchip_memory_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_001:sink_endofpacket
	wire         onchip_memory_s1_translator_avalon_universal_slave_0_agent_rp_valid;                               // onchip_memory_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_001:sink_valid
	wire         onchip_memory_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket;                       // onchip_memory_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_001:sink_startofpacket
	wire  [75:0] onchip_memory_s1_translator_avalon_universal_slave_0_agent_rp_data;                                // onchip_memory_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_001:sink_data
	wire         onchip_memory_s1_translator_avalon_universal_slave_0_agent_rp_ready;                               // id_router_001:sink_ready -> onchip_memory_s1_translator_avalon_universal_slave_0_agent:rp_ready
	wire         jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket;              // jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_002:sink_endofpacket
	wire         jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_valid;                    // jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_002:sink_valid
	wire         jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket;            // jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_002:sink_startofpacket
	wire  [75:0] jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_data;                     // jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rp_data -> id_router_002:sink_data
	wire         jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_ready;                    // id_router_002:sink_ready -> jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rp_ready
	wire         sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket;                 // sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_003:sink_endofpacket
	wire         sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent_rp_valid;                       // sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_003:sink_valid
	wire         sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket;               // sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_003:sink_startofpacket
	wire  [75:0] sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent_rp_data;                        // sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent:rp_data -> id_router_003:sink_data
	wire         sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent_rp_ready;                       // id_router_003:sink_ready -> sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent:rp_ready
	wire         pio_ledg_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket;                              // pio_LEDG_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_004:sink_endofpacket
	wire         pio_ledg_s1_translator_avalon_universal_slave_0_agent_rp_valid;                                    // pio_LEDG_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_004:sink_valid
	wire         pio_ledg_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket;                            // pio_LEDG_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_004:sink_startofpacket
	wire  [75:0] pio_ledg_s1_translator_avalon_universal_slave_0_agent_rp_data;                                     // pio_LEDG_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_004:sink_data
	wire         pio_ledg_s1_translator_avalon_universal_slave_0_agent_rp_ready;                                    // id_router_004:sink_ready -> pio_LEDG_s1_translator_avalon_universal_slave_0_agent:rp_ready
	wire         pio_ledr_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket;                              // pio_LEDR_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_005:sink_endofpacket
	wire         pio_ledr_s1_translator_avalon_universal_slave_0_agent_rp_valid;                                    // pio_LEDR_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_005:sink_valid
	wire         pio_ledr_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket;                            // pio_LEDR_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_005:sink_startofpacket
	wire  [75:0] pio_ledr_s1_translator_avalon_universal_slave_0_agent_rp_data;                                     // pio_LEDR_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_005:sink_data
	wire         pio_ledr_s1_translator_avalon_universal_slave_0_agent_rp_ready;                                    // id_router_005:sink_ready -> pio_LEDR_s1_translator_avalon_universal_slave_0_agent:rp_ready
	wire         pio_sw_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket;                                // pio_SW_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_006:sink_endofpacket
	wire         pio_sw_s1_translator_avalon_universal_slave_0_agent_rp_valid;                                      // pio_SW_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_006:sink_valid
	wire         pio_sw_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket;                              // pio_SW_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_006:sink_startofpacket
	wire  [75:0] pio_sw_s1_translator_avalon_universal_slave_0_agent_rp_data;                                       // pio_SW_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_006:sink_data
	wire         pio_sw_s1_translator_avalon_universal_slave_0_agent_rp_ready;                                      // id_router_006:sink_ready -> pio_SW_s1_translator_avalon_universal_slave_0_agent:rp_ready
	wire         pio_button_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket;                            // pio_Button_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_007:sink_endofpacket
	wire         pio_button_s1_translator_avalon_universal_slave_0_agent_rp_valid;                                  // pio_Button_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_007:sink_valid
	wire         pio_button_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket;                          // pio_Button_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_007:sink_startofpacket
	wire  [75:0] pio_button_s1_translator_avalon_universal_slave_0_agent_rp_data;                                   // pio_Button_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_007:sink_data
	wire         pio_button_s1_translator_avalon_universal_slave_0_agent_rp_ready;                                  // id_router_007:sink_ready -> pio_Button_s1_translator_avalon_universal_slave_0_agent:rp_ready
	wire         lcd_control_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket;                        // lcd_control_slave_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_008:sink_endofpacket
	wire         lcd_control_slave_translator_avalon_universal_slave_0_agent_rp_valid;                              // lcd_control_slave_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_008:sink_valid
	wire         lcd_control_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket;                      // lcd_control_slave_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_008:sink_startofpacket
	wire  [75:0] lcd_control_slave_translator_avalon_universal_slave_0_agent_rp_data;                               // lcd_control_slave_translator_avalon_universal_slave_0_agent:rp_data -> id_router_008:sink_data
	wire         lcd_control_slave_translator_avalon_universal_slave_0_agent_rp_ready;                              // id_router_008:sink_ready -> lcd_control_slave_translator_avalon_universal_slave_0_agent:rp_ready
	wire         uart_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket;                                  // uart_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_009:sink_endofpacket
	wire         uart_s1_translator_avalon_universal_slave_0_agent_rp_valid;                                        // uart_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_009:sink_valid
	wire         uart_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket;                                // uart_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_009:sink_startofpacket
	wire  [75:0] uart_s1_translator_avalon_universal_slave_0_agent_rp_data;                                         // uart_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_009:sink_data
	wire         uart_s1_translator_avalon_universal_slave_0_agent_rp_ready;                                        // id_router_009:sink_ready -> uart_s1_translator_avalon_universal_slave_0_agent:rp_ready
	wire         timer_0_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket;                               // timer_0_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_010:sink_endofpacket
	wire         timer_0_s1_translator_avalon_universal_slave_0_agent_rp_valid;                                     // timer_0_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_010:sink_valid
	wire         timer_0_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket;                             // timer_0_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_010:sink_startofpacket
	wire  [75:0] timer_0_s1_translator_avalon_universal_slave_0_agent_rp_data;                                      // timer_0_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_010:sink_data
	wire         timer_0_s1_translator_avalon_universal_slave_0_agent_rp_ready;                                     // id_router_010:sink_ready -> timer_0_s1_translator_avalon_universal_slave_0_agent:rp_ready
	wire         pio_data_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket;                              // pio_Data_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_011:sink_endofpacket
	wire         pio_data_s1_translator_avalon_universal_slave_0_agent_rp_valid;                                    // pio_Data_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_011:sink_valid
	wire         pio_data_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket;                            // pio_Data_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_011:sink_startofpacket
	wire  [75:0] pio_data_s1_translator_avalon_universal_slave_0_agent_rp_data;                                     // pio_Data_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_011:sink_data
	wire         pio_data_s1_translator_avalon_universal_slave_0_agent_rp_ready;                                    // id_router_011:sink_ready -> pio_Data_s1_translator_avalon_universal_slave_0_agent:rp_ready
	wire         pio_rdydata_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket;                           // pio_RdyData_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_012:sink_endofpacket
	wire         pio_rdydata_s1_translator_avalon_universal_slave_0_agent_rp_valid;                                 // pio_RdyData_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_012:sink_valid
	wire         pio_rdydata_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket;                         // pio_RdyData_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_012:sink_startofpacket
	wire  [75:0] pio_rdydata_s1_translator_avalon_universal_slave_0_agent_rp_data;                                  // pio_RdyData_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_012:sink_data
	wire         pio_rdydata_s1_translator_avalon_universal_slave_0_agent_rp_ready;                                 // id_router_012:sink_ready -> pio_RdyData_s1_translator_avalon_universal_slave_0_agent:rp_ready
	wire         pio_dataread_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket;                          // pio_DataRead_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_013:sink_endofpacket
	wire         pio_dataread_s1_translator_avalon_universal_slave_0_agent_rp_valid;                                // pio_DataRead_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_013:sink_valid
	wire         pio_dataread_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket;                        // pio_DataRead_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_013:sink_startofpacket
	wire  [75:0] pio_dataread_s1_translator_avalon_universal_slave_0_agent_rp_data;                                 // pio_DataRead_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_013:sink_data
	wire         pio_dataread_s1_translator_avalon_universal_slave_0_agent_rp_ready;                                // id_router_013:sink_ready -> pio_DataRead_s1_translator_avalon_universal_slave_0_agent:rp_ready
	wire         addr_router_src_endofpacket;                                                                       // addr_router:src_endofpacket -> limiter:cmd_sink_endofpacket
	wire         addr_router_src_valid;                                                                             // addr_router:src_valid -> limiter:cmd_sink_valid
	wire         addr_router_src_startofpacket;                                                                     // addr_router:src_startofpacket -> limiter:cmd_sink_startofpacket
	wire  [75:0] addr_router_src_data;                                                                              // addr_router:src_data -> limiter:cmd_sink_data
	wire  [13:0] addr_router_src_channel;                                                                           // addr_router:src_channel -> limiter:cmd_sink_channel
	wire         addr_router_src_ready;                                                                             // limiter:cmd_sink_ready -> addr_router:src_ready
	wire         limiter_rsp_src_endofpacket;                                                                       // limiter:rsp_src_endofpacket -> nios2_qsys_instruction_master_translator_avalon_universal_master_0_agent:rp_endofpacket
	wire         limiter_rsp_src_valid;                                                                             // limiter:rsp_src_valid -> nios2_qsys_instruction_master_translator_avalon_universal_master_0_agent:rp_valid
	wire         limiter_rsp_src_startofpacket;                                                                     // limiter:rsp_src_startofpacket -> nios2_qsys_instruction_master_translator_avalon_universal_master_0_agent:rp_startofpacket
	wire  [75:0] limiter_rsp_src_data;                                                                              // limiter:rsp_src_data -> nios2_qsys_instruction_master_translator_avalon_universal_master_0_agent:rp_data
	wire  [13:0] limiter_rsp_src_channel;                                                                           // limiter:rsp_src_channel -> nios2_qsys_instruction_master_translator_avalon_universal_master_0_agent:rp_channel
	wire         limiter_rsp_src_ready;                                                                             // nios2_qsys_instruction_master_translator_avalon_universal_master_0_agent:rp_ready -> limiter:rsp_src_ready
	wire         addr_router_001_src_endofpacket;                                                                   // addr_router_001:src_endofpacket -> limiter_001:cmd_sink_endofpacket
	wire         addr_router_001_src_valid;                                                                         // addr_router_001:src_valid -> limiter_001:cmd_sink_valid
	wire         addr_router_001_src_startofpacket;                                                                 // addr_router_001:src_startofpacket -> limiter_001:cmd_sink_startofpacket
	wire  [75:0] addr_router_001_src_data;                                                                          // addr_router_001:src_data -> limiter_001:cmd_sink_data
	wire  [13:0] addr_router_001_src_channel;                                                                       // addr_router_001:src_channel -> limiter_001:cmd_sink_channel
	wire         addr_router_001_src_ready;                                                                         // limiter_001:cmd_sink_ready -> addr_router_001:src_ready
	wire         limiter_001_rsp_src_endofpacket;                                                                   // limiter_001:rsp_src_endofpacket -> nios2_qsys_data_master_translator_avalon_universal_master_0_agent:rp_endofpacket
	wire         limiter_001_rsp_src_valid;                                                                         // limiter_001:rsp_src_valid -> nios2_qsys_data_master_translator_avalon_universal_master_0_agent:rp_valid
	wire         limiter_001_rsp_src_startofpacket;                                                                 // limiter_001:rsp_src_startofpacket -> nios2_qsys_data_master_translator_avalon_universal_master_0_agent:rp_startofpacket
	wire  [75:0] limiter_001_rsp_src_data;                                                                          // limiter_001:rsp_src_data -> nios2_qsys_data_master_translator_avalon_universal_master_0_agent:rp_data
	wire  [13:0] limiter_001_rsp_src_channel;                                                                       // limiter_001:rsp_src_channel -> nios2_qsys_data_master_translator_avalon_universal_master_0_agent:rp_channel
	wire         limiter_001_rsp_src_ready;                                                                         // nios2_qsys_data_master_translator_avalon_universal_master_0_agent:rp_ready -> limiter_001:rsp_src_ready
	wire         rst_controller_reset_out_reset;                                                                    // rst_controller:reset_out -> [addr_router:reset, addr_router_001:reset, cmd_xbar_demux:reset, cmd_xbar_demux_001:reset, cmd_xbar_mux:reset, cmd_xbar_mux_001:reset, id_router:reset, id_router_001:reset, id_router_002:reset, id_router_003:reset, id_router_004:reset, id_router_005:reset, id_router_006:reset, id_router_007:reset, id_router_008:reset, id_router_009:reset, id_router_010:reset, id_router_011:reset, id_router_012:reset, id_router_013:reset, irq_mapper:reset, jtag_uart:rst_n, jtag_uart_avalon_jtag_slave_translator:reset, jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:reset, jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, lcd:reset_n, lcd_control_slave_translator:reset, lcd_control_slave_translator_avalon_universal_slave_0_agent:reset, lcd_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, limiter:reset, limiter_001:reset, nios2_qsys:reset_n, nios2_qsys_data_master_translator:reset, nios2_qsys_data_master_translator_avalon_universal_master_0_agent:reset, nios2_qsys_instruction_master_translator:reset, nios2_qsys_instruction_master_translator_avalon_universal_master_0_agent:reset, nios2_qsys_jtag_debug_module_translator:reset, nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent:reset, nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, onchip_memory:reset, onchip_memory_s1_translator:reset, onchip_memory_s1_translator_avalon_universal_slave_0_agent:reset, onchip_memory_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, pio_Button:reset_n, pio_Button_s1_translator:reset, pio_Button_s1_translator_avalon_universal_slave_0_agent:reset, pio_Button_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, pio_Data:reset_n, pio_DataRead:reset_n, pio_DataRead_s1_translator:reset, pio_DataRead_s1_translator_avalon_universal_slave_0_agent:reset, pio_DataRead_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, pio_Data_s1_translator:reset, pio_Data_s1_translator_avalon_universal_slave_0_agent:reset, pio_Data_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, pio_LEDG:reset_n, pio_LEDG_s1_translator:reset, pio_LEDG_s1_translator_avalon_universal_slave_0_agent:reset, pio_LEDG_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, pio_LEDR:reset_n, pio_LEDR_s1_translator:reset, pio_LEDR_s1_translator_avalon_universal_slave_0_agent:reset, pio_LEDR_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, pio_RdyData:reset_n, pio_RdyData_s1_translator:reset, pio_RdyData_s1_translator_avalon_universal_slave_0_agent:reset, pio_RdyData_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, pio_SW:reset_n, pio_SW_s1_translator:reset, pio_SW_s1_translator_avalon_universal_slave_0_agent:reset, pio_SW_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, rsp_xbar_demux:reset, rsp_xbar_demux_001:reset, rsp_xbar_demux_002:reset, rsp_xbar_demux_003:reset, rsp_xbar_demux_004:reset, rsp_xbar_demux_005:reset, rsp_xbar_demux_006:reset, rsp_xbar_demux_007:reset, rsp_xbar_demux_008:reset, rsp_xbar_demux_009:reset, rsp_xbar_demux_010:reset, rsp_xbar_demux_011:reset, rsp_xbar_demux_012:reset, rsp_xbar_demux_013:reset, rsp_xbar_mux:reset, rsp_xbar_mux_001:reset, sysid_qsys:reset_n, sysid_qsys_control_slave_translator:reset, sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent:reset, sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, timer_0:reset_n, timer_0_s1_translator:reset, timer_0_s1_translator_avalon_universal_slave_0_agent:reset, timer_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, uart:reset_n, uart_s1_translator:reset, uart_s1_translator_avalon_universal_slave_0_agent:reset, uart_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset]
	wire         cmd_xbar_demux_src0_endofpacket;                                                                   // cmd_xbar_demux:src0_endofpacket -> cmd_xbar_mux:sink0_endofpacket
	wire         cmd_xbar_demux_src0_valid;                                                                         // cmd_xbar_demux:src0_valid -> cmd_xbar_mux:sink0_valid
	wire         cmd_xbar_demux_src0_startofpacket;                                                                 // cmd_xbar_demux:src0_startofpacket -> cmd_xbar_mux:sink0_startofpacket
	wire  [75:0] cmd_xbar_demux_src0_data;                                                                          // cmd_xbar_demux:src0_data -> cmd_xbar_mux:sink0_data
	wire  [13:0] cmd_xbar_demux_src0_channel;                                                                       // cmd_xbar_demux:src0_channel -> cmd_xbar_mux:sink0_channel
	wire         cmd_xbar_demux_src0_ready;                                                                         // cmd_xbar_mux:sink0_ready -> cmd_xbar_demux:src0_ready
	wire         cmd_xbar_demux_src1_endofpacket;                                                                   // cmd_xbar_demux:src1_endofpacket -> cmd_xbar_mux_001:sink0_endofpacket
	wire         cmd_xbar_demux_src1_valid;                                                                         // cmd_xbar_demux:src1_valid -> cmd_xbar_mux_001:sink0_valid
	wire         cmd_xbar_demux_src1_startofpacket;                                                                 // cmd_xbar_demux:src1_startofpacket -> cmd_xbar_mux_001:sink0_startofpacket
	wire  [75:0] cmd_xbar_demux_src1_data;                                                                          // cmd_xbar_demux:src1_data -> cmd_xbar_mux_001:sink0_data
	wire  [13:0] cmd_xbar_demux_src1_channel;                                                                       // cmd_xbar_demux:src1_channel -> cmd_xbar_mux_001:sink0_channel
	wire         cmd_xbar_demux_src1_ready;                                                                         // cmd_xbar_mux_001:sink0_ready -> cmd_xbar_demux:src1_ready
	wire         cmd_xbar_demux_001_src0_endofpacket;                                                               // cmd_xbar_demux_001:src0_endofpacket -> cmd_xbar_mux:sink1_endofpacket
	wire         cmd_xbar_demux_001_src0_valid;                                                                     // cmd_xbar_demux_001:src0_valid -> cmd_xbar_mux:sink1_valid
	wire         cmd_xbar_demux_001_src0_startofpacket;                                                             // cmd_xbar_demux_001:src0_startofpacket -> cmd_xbar_mux:sink1_startofpacket
	wire  [75:0] cmd_xbar_demux_001_src0_data;                                                                      // cmd_xbar_demux_001:src0_data -> cmd_xbar_mux:sink1_data
	wire  [13:0] cmd_xbar_demux_001_src0_channel;                                                                   // cmd_xbar_demux_001:src0_channel -> cmd_xbar_mux:sink1_channel
	wire         cmd_xbar_demux_001_src0_ready;                                                                     // cmd_xbar_mux:sink1_ready -> cmd_xbar_demux_001:src0_ready
	wire         cmd_xbar_demux_001_src1_endofpacket;                                                               // cmd_xbar_demux_001:src1_endofpacket -> cmd_xbar_mux_001:sink1_endofpacket
	wire         cmd_xbar_demux_001_src1_valid;                                                                     // cmd_xbar_demux_001:src1_valid -> cmd_xbar_mux_001:sink1_valid
	wire         cmd_xbar_demux_001_src1_startofpacket;                                                             // cmd_xbar_demux_001:src1_startofpacket -> cmd_xbar_mux_001:sink1_startofpacket
	wire  [75:0] cmd_xbar_demux_001_src1_data;                                                                      // cmd_xbar_demux_001:src1_data -> cmd_xbar_mux_001:sink1_data
	wire  [13:0] cmd_xbar_demux_001_src1_channel;                                                                   // cmd_xbar_demux_001:src1_channel -> cmd_xbar_mux_001:sink1_channel
	wire         cmd_xbar_demux_001_src1_ready;                                                                     // cmd_xbar_mux_001:sink1_ready -> cmd_xbar_demux_001:src1_ready
	wire         cmd_xbar_demux_001_src2_endofpacket;                                                               // cmd_xbar_demux_001:src2_endofpacket -> jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire         cmd_xbar_demux_001_src2_valid;                                                                     // cmd_xbar_demux_001:src2_valid -> jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:cp_valid
	wire         cmd_xbar_demux_001_src2_startofpacket;                                                             // cmd_xbar_demux_001:src2_startofpacket -> jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [75:0] cmd_xbar_demux_001_src2_data;                                                                      // cmd_xbar_demux_001:src2_data -> jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:cp_data
	wire  [13:0] cmd_xbar_demux_001_src2_channel;                                                                   // cmd_xbar_demux_001:src2_channel -> jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:cp_channel
	wire         cmd_xbar_demux_001_src3_endofpacket;                                                               // cmd_xbar_demux_001:src3_endofpacket -> sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire         cmd_xbar_demux_001_src3_valid;                                                                     // cmd_xbar_demux_001:src3_valid -> sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent:cp_valid
	wire         cmd_xbar_demux_001_src3_startofpacket;                                                             // cmd_xbar_demux_001:src3_startofpacket -> sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [75:0] cmd_xbar_demux_001_src3_data;                                                                      // cmd_xbar_demux_001:src3_data -> sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent:cp_data
	wire  [13:0] cmd_xbar_demux_001_src3_channel;                                                                   // cmd_xbar_demux_001:src3_channel -> sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent:cp_channel
	wire         cmd_xbar_demux_001_src4_endofpacket;                                                               // cmd_xbar_demux_001:src4_endofpacket -> pio_LEDG_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire         cmd_xbar_demux_001_src4_valid;                                                                     // cmd_xbar_demux_001:src4_valid -> pio_LEDG_s1_translator_avalon_universal_slave_0_agent:cp_valid
	wire         cmd_xbar_demux_001_src4_startofpacket;                                                             // cmd_xbar_demux_001:src4_startofpacket -> pio_LEDG_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [75:0] cmd_xbar_demux_001_src4_data;                                                                      // cmd_xbar_demux_001:src4_data -> pio_LEDG_s1_translator_avalon_universal_slave_0_agent:cp_data
	wire  [13:0] cmd_xbar_demux_001_src4_channel;                                                                   // cmd_xbar_demux_001:src4_channel -> pio_LEDG_s1_translator_avalon_universal_slave_0_agent:cp_channel
	wire         cmd_xbar_demux_001_src5_endofpacket;                                                               // cmd_xbar_demux_001:src5_endofpacket -> pio_LEDR_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire         cmd_xbar_demux_001_src5_valid;                                                                     // cmd_xbar_demux_001:src5_valid -> pio_LEDR_s1_translator_avalon_universal_slave_0_agent:cp_valid
	wire         cmd_xbar_demux_001_src5_startofpacket;                                                             // cmd_xbar_demux_001:src5_startofpacket -> pio_LEDR_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [75:0] cmd_xbar_demux_001_src5_data;                                                                      // cmd_xbar_demux_001:src5_data -> pio_LEDR_s1_translator_avalon_universal_slave_0_agent:cp_data
	wire  [13:0] cmd_xbar_demux_001_src5_channel;                                                                   // cmd_xbar_demux_001:src5_channel -> pio_LEDR_s1_translator_avalon_universal_slave_0_agent:cp_channel
	wire         cmd_xbar_demux_001_src6_endofpacket;                                                               // cmd_xbar_demux_001:src6_endofpacket -> pio_SW_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire         cmd_xbar_demux_001_src6_valid;                                                                     // cmd_xbar_demux_001:src6_valid -> pio_SW_s1_translator_avalon_universal_slave_0_agent:cp_valid
	wire         cmd_xbar_demux_001_src6_startofpacket;                                                             // cmd_xbar_demux_001:src6_startofpacket -> pio_SW_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [75:0] cmd_xbar_demux_001_src6_data;                                                                      // cmd_xbar_demux_001:src6_data -> pio_SW_s1_translator_avalon_universal_slave_0_agent:cp_data
	wire  [13:0] cmd_xbar_demux_001_src6_channel;                                                                   // cmd_xbar_demux_001:src6_channel -> pio_SW_s1_translator_avalon_universal_slave_0_agent:cp_channel
	wire         cmd_xbar_demux_001_src7_endofpacket;                                                               // cmd_xbar_demux_001:src7_endofpacket -> pio_Button_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire         cmd_xbar_demux_001_src7_valid;                                                                     // cmd_xbar_demux_001:src7_valid -> pio_Button_s1_translator_avalon_universal_slave_0_agent:cp_valid
	wire         cmd_xbar_demux_001_src7_startofpacket;                                                             // cmd_xbar_demux_001:src7_startofpacket -> pio_Button_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [75:0] cmd_xbar_demux_001_src7_data;                                                                      // cmd_xbar_demux_001:src7_data -> pio_Button_s1_translator_avalon_universal_slave_0_agent:cp_data
	wire  [13:0] cmd_xbar_demux_001_src7_channel;                                                                   // cmd_xbar_demux_001:src7_channel -> pio_Button_s1_translator_avalon_universal_slave_0_agent:cp_channel
	wire         cmd_xbar_demux_001_src8_endofpacket;                                                               // cmd_xbar_demux_001:src8_endofpacket -> lcd_control_slave_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire         cmd_xbar_demux_001_src8_valid;                                                                     // cmd_xbar_demux_001:src8_valid -> lcd_control_slave_translator_avalon_universal_slave_0_agent:cp_valid
	wire         cmd_xbar_demux_001_src8_startofpacket;                                                             // cmd_xbar_demux_001:src8_startofpacket -> lcd_control_slave_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [75:0] cmd_xbar_demux_001_src8_data;                                                                      // cmd_xbar_demux_001:src8_data -> lcd_control_slave_translator_avalon_universal_slave_0_agent:cp_data
	wire  [13:0] cmd_xbar_demux_001_src8_channel;                                                                   // cmd_xbar_demux_001:src8_channel -> lcd_control_slave_translator_avalon_universal_slave_0_agent:cp_channel
	wire         cmd_xbar_demux_001_src9_endofpacket;                                                               // cmd_xbar_demux_001:src9_endofpacket -> uart_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire         cmd_xbar_demux_001_src9_valid;                                                                     // cmd_xbar_demux_001:src9_valid -> uart_s1_translator_avalon_universal_slave_0_agent:cp_valid
	wire         cmd_xbar_demux_001_src9_startofpacket;                                                             // cmd_xbar_demux_001:src9_startofpacket -> uart_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [75:0] cmd_xbar_demux_001_src9_data;                                                                      // cmd_xbar_demux_001:src9_data -> uart_s1_translator_avalon_universal_slave_0_agent:cp_data
	wire  [13:0] cmd_xbar_demux_001_src9_channel;                                                                   // cmd_xbar_demux_001:src9_channel -> uart_s1_translator_avalon_universal_slave_0_agent:cp_channel
	wire         cmd_xbar_demux_001_src10_endofpacket;                                                              // cmd_xbar_demux_001:src10_endofpacket -> timer_0_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire         cmd_xbar_demux_001_src10_valid;                                                                    // cmd_xbar_demux_001:src10_valid -> timer_0_s1_translator_avalon_universal_slave_0_agent:cp_valid
	wire         cmd_xbar_demux_001_src10_startofpacket;                                                            // cmd_xbar_demux_001:src10_startofpacket -> timer_0_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [75:0] cmd_xbar_demux_001_src10_data;                                                                     // cmd_xbar_demux_001:src10_data -> timer_0_s1_translator_avalon_universal_slave_0_agent:cp_data
	wire  [13:0] cmd_xbar_demux_001_src10_channel;                                                                  // cmd_xbar_demux_001:src10_channel -> timer_0_s1_translator_avalon_universal_slave_0_agent:cp_channel
	wire         cmd_xbar_demux_001_src11_endofpacket;                                                              // cmd_xbar_demux_001:src11_endofpacket -> pio_Data_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire         cmd_xbar_demux_001_src11_valid;                                                                    // cmd_xbar_demux_001:src11_valid -> pio_Data_s1_translator_avalon_universal_slave_0_agent:cp_valid
	wire         cmd_xbar_demux_001_src11_startofpacket;                                                            // cmd_xbar_demux_001:src11_startofpacket -> pio_Data_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [75:0] cmd_xbar_demux_001_src11_data;                                                                     // cmd_xbar_demux_001:src11_data -> pio_Data_s1_translator_avalon_universal_slave_0_agent:cp_data
	wire  [13:0] cmd_xbar_demux_001_src11_channel;                                                                  // cmd_xbar_demux_001:src11_channel -> pio_Data_s1_translator_avalon_universal_slave_0_agent:cp_channel
	wire         cmd_xbar_demux_001_src12_endofpacket;                                                              // cmd_xbar_demux_001:src12_endofpacket -> pio_RdyData_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire         cmd_xbar_demux_001_src12_valid;                                                                    // cmd_xbar_demux_001:src12_valid -> pio_RdyData_s1_translator_avalon_universal_slave_0_agent:cp_valid
	wire         cmd_xbar_demux_001_src12_startofpacket;                                                            // cmd_xbar_demux_001:src12_startofpacket -> pio_RdyData_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [75:0] cmd_xbar_demux_001_src12_data;                                                                     // cmd_xbar_demux_001:src12_data -> pio_RdyData_s1_translator_avalon_universal_slave_0_agent:cp_data
	wire  [13:0] cmd_xbar_demux_001_src12_channel;                                                                  // cmd_xbar_demux_001:src12_channel -> pio_RdyData_s1_translator_avalon_universal_slave_0_agent:cp_channel
	wire         cmd_xbar_demux_001_src13_endofpacket;                                                              // cmd_xbar_demux_001:src13_endofpacket -> pio_DataRead_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire         cmd_xbar_demux_001_src13_valid;                                                                    // cmd_xbar_demux_001:src13_valid -> pio_DataRead_s1_translator_avalon_universal_slave_0_agent:cp_valid
	wire         cmd_xbar_demux_001_src13_startofpacket;                                                            // cmd_xbar_demux_001:src13_startofpacket -> pio_DataRead_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [75:0] cmd_xbar_demux_001_src13_data;                                                                     // cmd_xbar_demux_001:src13_data -> pio_DataRead_s1_translator_avalon_universal_slave_0_agent:cp_data
	wire  [13:0] cmd_xbar_demux_001_src13_channel;                                                                  // cmd_xbar_demux_001:src13_channel -> pio_DataRead_s1_translator_avalon_universal_slave_0_agent:cp_channel
	wire         rsp_xbar_demux_src0_endofpacket;                                                                   // rsp_xbar_demux:src0_endofpacket -> rsp_xbar_mux:sink0_endofpacket
	wire         rsp_xbar_demux_src0_valid;                                                                         // rsp_xbar_demux:src0_valid -> rsp_xbar_mux:sink0_valid
	wire         rsp_xbar_demux_src0_startofpacket;                                                                 // rsp_xbar_demux:src0_startofpacket -> rsp_xbar_mux:sink0_startofpacket
	wire  [75:0] rsp_xbar_demux_src0_data;                                                                          // rsp_xbar_demux:src0_data -> rsp_xbar_mux:sink0_data
	wire  [13:0] rsp_xbar_demux_src0_channel;                                                                       // rsp_xbar_demux:src0_channel -> rsp_xbar_mux:sink0_channel
	wire         rsp_xbar_demux_src0_ready;                                                                         // rsp_xbar_mux:sink0_ready -> rsp_xbar_demux:src0_ready
	wire         rsp_xbar_demux_src1_endofpacket;                                                                   // rsp_xbar_demux:src1_endofpacket -> rsp_xbar_mux_001:sink0_endofpacket
	wire         rsp_xbar_demux_src1_valid;                                                                         // rsp_xbar_demux:src1_valid -> rsp_xbar_mux_001:sink0_valid
	wire         rsp_xbar_demux_src1_startofpacket;                                                                 // rsp_xbar_demux:src1_startofpacket -> rsp_xbar_mux_001:sink0_startofpacket
	wire  [75:0] rsp_xbar_demux_src1_data;                                                                          // rsp_xbar_demux:src1_data -> rsp_xbar_mux_001:sink0_data
	wire  [13:0] rsp_xbar_demux_src1_channel;                                                                       // rsp_xbar_demux:src1_channel -> rsp_xbar_mux_001:sink0_channel
	wire         rsp_xbar_demux_src1_ready;                                                                         // rsp_xbar_mux_001:sink0_ready -> rsp_xbar_demux:src1_ready
	wire         rsp_xbar_demux_001_src0_endofpacket;                                                               // rsp_xbar_demux_001:src0_endofpacket -> rsp_xbar_mux:sink1_endofpacket
	wire         rsp_xbar_demux_001_src0_valid;                                                                     // rsp_xbar_demux_001:src0_valid -> rsp_xbar_mux:sink1_valid
	wire         rsp_xbar_demux_001_src0_startofpacket;                                                             // rsp_xbar_demux_001:src0_startofpacket -> rsp_xbar_mux:sink1_startofpacket
	wire  [75:0] rsp_xbar_demux_001_src0_data;                                                                      // rsp_xbar_demux_001:src0_data -> rsp_xbar_mux:sink1_data
	wire  [13:0] rsp_xbar_demux_001_src0_channel;                                                                   // rsp_xbar_demux_001:src0_channel -> rsp_xbar_mux:sink1_channel
	wire         rsp_xbar_demux_001_src0_ready;                                                                     // rsp_xbar_mux:sink1_ready -> rsp_xbar_demux_001:src0_ready
	wire         rsp_xbar_demux_001_src1_endofpacket;                                                               // rsp_xbar_demux_001:src1_endofpacket -> rsp_xbar_mux_001:sink1_endofpacket
	wire         rsp_xbar_demux_001_src1_valid;                                                                     // rsp_xbar_demux_001:src1_valid -> rsp_xbar_mux_001:sink1_valid
	wire         rsp_xbar_demux_001_src1_startofpacket;                                                             // rsp_xbar_demux_001:src1_startofpacket -> rsp_xbar_mux_001:sink1_startofpacket
	wire  [75:0] rsp_xbar_demux_001_src1_data;                                                                      // rsp_xbar_demux_001:src1_data -> rsp_xbar_mux_001:sink1_data
	wire  [13:0] rsp_xbar_demux_001_src1_channel;                                                                   // rsp_xbar_demux_001:src1_channel -> rsp_xbar_mux_001:sink1_channel
	wire         rsp_xbar_demux_001_src1_ready;                                                                     // rsp_xbar_mux_001:sink1_ready -> rsp_xbar_demux_001:src1_ready
	wire         rsp_xbar_demux_002_src0_endofpacket;                                                               // rsp_xbar_demux_002:src0_endofpacket -> rsp_xbar_mux_001:sink2_endofpacket
	wire         rsp_xbar_demux_002_src0_valid;                                                                     // rsp_xbar_demux_002:src0_valid -> rsp_xbar_mux_001:sink2_valid
	wire         rsp_xbar_demux_002_src0_startofpacket;                                                             // rsp_xbar_demux_002:src0_startofpacket -> rsp_xbar_mux_001:sink2_startofpacket
	wire  [75:0] rsp_xbar_demux_002_src0_data;                                                                      // rsp_xbar_demux_002:src0_data -> rsp_xbar_mux_001:sink2_data
	wire  [13:0] rsp_xbar_demux_002_src0_channel;                                                                   // rsp_xbar_demux_002:src0_channel -> rsp_xbar_mux_001:sink2_channel
	wire         rsp_xbar_demux_002_src0_ready;                                                                     // rsp_xbar_mux_001:sink2_ready -> rsp_xbar_demux_002:src0_ready
	wire         rsp_xbar_demux_003_src0_endofpacket;                                                               // rsp_xbar_demux_003:src0_endofpacket -> rsp_xbar_mux_001:sink3_endofpacket
	wire         rsp_xbar_demux_003_src0_valid;                                                                     // rsp_xbar_demux_003:src0_valid -> rsp_xbar_mux_001:sink3_valid
	wire         rsp_xbar_demux_003_src0_startofpacket;                                                             // rsp_xbar_demux_003:src0_startofpacket -> rsp_xbar_mux_001:sink3_startofpacket
	wire  [75:0] rsp_xbar_demux_003_src0_data;                                                                      // rsp_xbar_demux_003:src0_data -> rsp_xbar_mux_001:sink3_data
	wire  [13:0] rsp_xbar_demux_003_src0_channel;                                                                   // rsp_xbar_demux_003:src0_channel -> rsp_xbar_mux_001:sink3_channel
	wire         rsp_xbar_demux_003_src0_ready;                                                                     // rsp_xbar_mux_001:sink3_ready -> rsp_xbar_demux_003:src0_ready
	wire         rsp_xbar_demux_004_src0_endofpacket;                                                               // rsp_xbar_demux_004:src0_endofpacket -> rsp_xbar_mux_001:sink4_endofpacket
	wire         rsp_xbar_demux_004_src0_valid;                                                                     // rsp_xbar_demux_004:src0_valid -> rsp_xbar_mux_001:sink4_valid
	wire         rsp_xbar_demux_004_src0_startofpacket;                                                             // rsp_xbar_demux_004:src0_startofpacket -> rsp_xbar_mux_001:sink4_startofpacket
	wire  [75:0] rsp_xbar_demux_004_src0_data;                                                                      // rsp_xbar_demux_004:src0_data -> rsp_xbar_mux_001:sink4_data
	wire  [13:0] rsp_xbar_demux_004_src0_channel;                                                                   // rsp_xbar_demux_004:src0_channel -> rsp_xbar_mux_001:sink4_channel
	wire         rsp_xbar_demux_004_src0_ready;                                                                     // rsp_xbar_mux_001:sink4_ready -> rsp_xbar_demux_004:src0_ready
	wire         rsp_xbar_demux_005_src0_endofpacket;                                                               // rsp_xbar_demux_005:src0_endofpacket -> rsp_xbar_mux_001:sink5_endofpacket
	wire         rsp_xbar_demux_005_src0_valid;                                                                     // rsp_xbar_demux_005:src0_valid -> rsp_xbar_mux_001:sink5_valid
	wire         rsp_xbar_demux_005_src0_startofpacket;                                                             // rsp_xbar_demux_005:src0_startofpacket -> rsp_xbar_mux_001:sink5_startofpacket
	wire  [75:0] rsp_xbar_demux_005_src0_data;                                                                      // rsp_xbar_demux_005:src0_data -> rsp_xbar_mux_001:sink5_data
	wire  [13:0] rsp_xbar_demux_005_src0_channel;                                                                   // rsp_xbar_demux_005:src0_channel -> rsp_xbar_mux_001:sink5_channel
	wire         rsp_xbar_demux_005_src0_ready;                                                                     // rsp_xbar_mux_001:sink5_ready -> rsp_xbar_demux_005:src0_ready
	wire         rsp_xbar_demux_006_src0_endofpacket;                                                               // rsp_xbar_demux_006:src0_endofpacket -> rsp_xbar_mux_001:sink6_endofpacket
	wire         rsp_xbar_demux_006_src0_valid;                                                                     // rsp_xbar_demux_006:src0_valid -> rsp_xbar_mux_001:sink6_valid
	wire         rsp_xbar_demux_006_src0_startofpacket;                                                             // rsp_xbar_demux_006:src0_startofpacket -> rsp_xbar_mux_001:sink6_startofpacket
	wire  [75:0] rsp_xbar_demux_006_src0_data;                                                                      // rsp_xbar_demux_006:src0_data -> rsp_xbar_mux_001:sink6_data
	wire  [13:0] rsp_xbar_demux_006_src0_channel;                                                                   // rsp_xbar_demux_006:src0_channel -> rsp_xbar_mux_001:sink6_channel
	wire         rsp_xbar_demux_006_src0_ready;                                                                     // rsp_xbar_mux_001:sink6_ready -> rsp_xbar_demux_006:src0_ready
	wire         rsp_xbar_demux_007_src0_endofpacket;                                                               // rsp_xbar_demux_007:src0_endofpacket -> rsp_xbar_mux_001:sink7_endofpacket
	wire         rsp_xbar_demux_007_src0_valid;                                                                     // rsp_xbar_demux_007:src0_valid -> rsp_xbar_mux_001:sink7_valid
	wire         rsp_xbar_demux_007_src0_startofpacket;                                                             // rsp_xbar_demux_007:src0_startofpacket -> rsp_xbar_mux_001:sink7_startofpacket
	wire  [75:0] rsp_xbar_demux_007_src0_data;                                                                      // rsp_xbar_demux_007:src0_data -> rsp_xbar_mux_001:sink7_data
	wire  [13:0] rsp_xbar_demux_007_src0_channel;                                                                   // rsp_xbar_demux_007:src0_channel -> rsp_xbar_mux_001:sink7_channel
	wire         rsp_xbar_demux_007_src0_ready;                                                                     // rsp_xbar_mux_001:sink7_ready -> rsp_xbar_demux_007:src0_ready
	wire         rsp_xbar_demux_008_src0_endofpacket;                                                               // rsp_xbar_demux_008:src0_endofpacket -> rsp_xbar_mux_001:sink8_endofpacket
	wire         rsp_xbar_demux_008_src0_valid;                                                                     // rsp_xbar_demux_008:src0_valid -> rsp_xbar_mux_001:sink8_valid
	wire         rsp_xbar_demux_008_src0_startofpacket;                                                             // rsp_xbar_demux_008:src0_startofpacket -> rsp_xbar_mux_001:sink8_startofpacket
	wire  [75:0] rsp_xbar_demux_008_src0_data;                                                                      // rsp_xbar_demux_008:src0_data -> rsp_xbar_mux_001:sink8_data
	wire  [13:0] rsp_xbar_demux_008_src0_channel;                                                                   // rsp_xbar_demux_008:src0_channel -> rsp_xbar_mux_001:sink8_channel
	wire         rsp_xbar_demux_008_src0_ready;                                                                     // rsp_xbar_mux_001:sink8_ready -> rsp_xbar_demux_008:src0_ready
	wire         rsp_xbar_demux_009_src0_endofpacket;                                                               // rsp_xbar_demux_009:src0_endofpacket -> rsp_xbar_mux_001:sink9_endofpacket
	wire         rsp_xbar_demux_009_src0_valid;                                                                     // rsp_xbar_demux_009:src0_valid -> rsp_xbar_mux_001:sink9_valid
	wire         rsp_xbar_demux_009_src0_startofpacket;                                                             // rsp_xbar_demux_009:src0_startofpacket -> rsp_xbar_mux_001:sink9_startofpacket
	wire  [75:0] rsp_xbar_demux_009_src0_data;                                                                      // rsp_xbar_demux_009:src0_data -> rsp_xbar_mux_001:sink9_data
	wire  [13:0] rsp_xbar_demux_009_src0_channel;                                                                   // rsp_xbar_demux_009:src0_channel -> rsp_xbar_mux_001:sink9_channel
	wire         rsp_xbar_demux_009_src0_ready;                                                                     // rsp_xbar_mux_001:sink9_ready -> rsp_xbar_demux_009:src0_ready
	wire         rsp_xbar_demux_010_src0_endofpacket;                                                               // rsp_xbar_demux_010:src0_endofpacket -> rsp_xbar_mux_001:sink10_endofpacket
	wire         rsp_xbar_demux_010_src0_valid;                                                                     // rsp_xbar_demux_010:src0_valid -> rsp_xbar_mux_001:sink10_valid
	wire         rsp_xbar_demux_010_src0_startofpacket;                                                             // rsp_xbar_demux_010:src0_startofpacket -> rsp_xbar_mux_001:sink10_startofpacket
	wire  [75:0] rsp_xbar_demux_010_src0_data;                                                                      // rsp_xbar_demux_010:src0_data -> rsp_xbar_mux_001:sink10_data
	wire  [13:0] rsp_xbar_demux_010_src0_channel;                                                                   // rsp_xbar_demux_010:src0_channel -> rsp_xbar_mux_001:sink10_channel
	wire         rsp_xbar_demux_010_src0_ready;                                                                     // rsp_xbar_mux_001:sink10_ready -> rsp_xbar_demux_010:src0_ready
	wire         rsp_xbar_demux_011_src0_endofpacket;                                                               // rsp_xbar_demux_011:src0_endofpacket -> rsp_xbar_mux_001:sink11_endofpacket
	wire         rsp_xbar_demux_011_src0_valid;                                                                     // rsp_xbar_demux_011:src0_valid -> rsp_xbar_mux_001:sink11_valid
	wire         rsp_xbar_demux_011_src0_startofpacket;                                                             // rsp_xbar_demux_011:src0_startofpacket -> rsp_xbar_mux_001:sink11_startofpacket
	wire  [75:0] rsp_xbar_demux_011_src0_data;                                                                      // rsp_xbar_demux_011:src0_data -> rsp_xbar_mux_001:sink11_data
	wire  [13:0] rsp_xbar_demux_011_src0_channel;                                                                   // rsp_xbar_demux_011:src0_channel -> rsp_xbar_mux_001:sink11_channel
	wire         rsp_xbar_demux_011_src0_ready;                                                                     // rsp_xbar_mux_001:sink11_ready -> rsp_xbar_demux_011:src0_ready
	wire         rsp_xbar_demux_012_src0_endofpacket;                                                               // rsp_xbar_demux_012:src0_endofpacket -> rsp_xbar_mux_001:sink12_endofpacket
	wire         rsp_xbar_demux_012_src0_valid;                                                                     // rsp_xbar_demux_012:src0_valid -> rsp_xbar_mux_001:sink12_valid
	wire         rsp_xbar_demux_012_src0_startofpacket;                                                             // rsp_xbar_demux_012:src0_startofpacket -> rsp_xbar_mux_001:sink12_startofpacket
	wire  [75:0] rsp_xbar_demux_012_src0_data;                                                                      // rsp_xbar_demux_012:src0_data -> rsp_xbar_mux_001:sink12_data
	wire  [13:0] rsp_xbar_demux_012_src0_channel;                                                                   // rsp_xbar_demux_012:src0_channel -> rsp_xbar_mux_001:sink12_channel
	wire         rsp_xbar_demux_012_src0_ready;                                                                     // rsp_xbar_mux_001:sink12_ready -> rsp_xbar_demux_012:src0_ready
	wire         rsp_xbar_demux_013_src0_endofpacket;                                                               // rsp_xbar_demux_013:src0_endofpacket -> rsp_xbar_mux_001:sink13_endofpacket
	wire         rsp_xbar_demux_013_src0_valid;                                                                     // rsp_xbar_demux_013:src0_valid -> rsp_xbar_mux_001:sink13_valid
	wire         rsp_xbar_demux_013_src0_startofpacket;                                                             // rsp_xbar_demux_013:src0_startofpacket -> rsp_xbar_mux_001:sink13_startofpacket
	wire  [75:0] rsp_xbar_demux_013_src0_data;                                                                      // rsp_xbar_demux_013:src0_data -> rsp_xbar_mux_001:sink13_data
	wire  [13:0] rsp_xbar_demux_013_src0_channel;                                                                   // rsp_xbar_demux_013:src0_channel -> rsp_xbar_mux_001:sink13_channel
	wire         rsp_xbar_demux_013_src0_ready;                                                                     // rsp_xbar_mux_001:sink13_ready -> rsp_xbar_demux_013:src0_ready
	wire         limiter_cmd_src_endofpacket;                                                                       // limiter:cmd_src_endofpacket -> cmd_xbar_demux:sink_endofpacket
	wire         limiter_cmd_src_startofpacket;                                                                     // limiter:cmd_src_startofpacket -> cmd_xbar_demux:sink_startofpacket
	wire  [75:0] limiter_cmd_src_data;                                                                              // limiter:cmd_src_data -> cmd_xbar_demux:sink_data
	wire  [13:0] limiter_cmd_src_channel;                                                                           // limiter:cmd_src_channel -> cmd_xbar_demux:sink_channel
	wire         limiter_cmd_src_ready;                                                                             // cmd_xbar_demux:sink_ready -> limiter:cmd_src_ready
	wire         rsp_xbar_mux_src_endofpacket;                                                                      // rsp_xbar_mux:src_endofpacket -> limiter:rsp_sink_endofpacket
	wire         rsp_xbar_mux_src_valid;                                                                            // rsp_xbar_mux:src_valid -> limiter:rsp_sink_valid
	wire         rsp_xbar_mux_src_startofpacket;                                                                    // rsp_xbar_mux:src_startofpacket -> limiter:rsp_sink_startofpacket
	wire  [75:0] rsp_xbar_mux_src_data;                                                                             // rsp_xbar_mux:src_data -> limiter:rsp_sink_data
	wire  [13:0] rsp_xbar_mux_src_channel;                                                                          // rsp_xbar_mux:src_channel -> limiter:rsp_sink_channel
	wire         rsp_xbar_mux_src_ready;                                                                            // limiter:rsp_sink_ready -> rsp_xbar_mux:src_ready
	wire         limiter_001_cmd_src_endofpacket;                                                                   // limiter_001:cmd_src_endofpacket -> cmd_xbar_demux_001:sink_endofpacket
	wire         limiter_001_cmd_src_startofpacket;                                                                 // limiter_001:cmd_src_startofpacket -> cmd_xbar_demux_001:sink_startofpacket
	wire  [75:0] limiter_001_cmd_src_data;                                                                          // limiter_001:cmd_src_data -> cmd_xbar_demux_001:sink_data
	wire  [13:0] limiter_001_cmd_src_channel;                                                                       // limiter_001:cmd_src_channel -> cmd_xbar_demux_001:sink_channel
	wire         limiter_001_cmd_src_ready;                                                                         // cmd_xbar_demux_001:sink_ready -> limiter_001:cmd_src_ready
	wire         rsp_xbar_mux_001_src_endofpacket;                                                                  // rsp_xbar_mux_001:src_endofpacket -> limiter_001:rsp_sink_endofpacket
	wire         rsp_xbar_mux_001_src_valid;                                                                        // rsp_xbar_mux_001:src_valid -> limiter_001:rsp_sink_valid
	wire         rsp_xbar_mux_001_src_startofpacket;                                                                // rsp_xbar_mux_001:src_startofpacket -> limiter_001:rsp_sink_startofpacket
	wire  [75:0] rsp_xbar_mux_001_src_data;                                                                         // rsp_xbar_mux_001:src_data -> limiter_001:rsp_sink_data
	wire  [13:0] rsp_xbar_mux_001_src_channel;                                                                      // rsp_xbar_mux_001:src_channel -> limiter_001:rsp_sink_channel
	wire         rsp_xbar_mux_001_src_ready;                                                                        // limiter_001:rsp_sink_ready -> rsp_xbar_mux_001:src_ready
	wire         cmd_xbar_mux_src_endofpacket;                                                                      // cmd_xbar_mux:src_endofpacket -> nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire         cmd_xbar_mux_src_valid;                                                                            // cmd_xbar_mux:src_valid -> nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent:cp_valid
	wire         cmd_xbar_mux_src_startofpacket;                                                                    // cmd_xbar_mux:src_startofpacket -> nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [75:0] cmd_xbar_mux_src_data;                                                                             // cmd_xbar_mux:src_data -> nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent:cp_data
	wire  [13:0] cmd_xbar_mux_src_channel;                                                                          // cmd_xbar_mux:src_channel -> nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent:cp_channel
	wire         cmd_xbar_mux_src_ready;                                                                            // nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_mux:src_ready
	wire         id_router_src_endofpacket;                                                                         // id_router:src_endofpacket -> rsp_xbar_demux:sink_endofpacket
	wire         id_router_src_valid;                                                                               // id_router:src_valid -> rsp_xbar_demux:sink_valid
	wire         id_router_src_startofpacket;                                                                       // id_router:src_startofpacket -> rsp_xbar_demux:sink_startofpacket
	wire  [75:0] id_router_src_data;                                                                                // id_router:src_data -> rsp_xbar_demux:sink_data
	wire  [13:0] id_router_src_channel;                                                                             // id_router:src_channel -> rsp_xbar_demux:sink_channel
	wire         id_router_src_ready;                                                                               // rsp_xbar_demux:sink_ready -> id_router:src_ready
	wire         cmd_xbar_mux_001_src_endofpacket;                                                                  // cmd_xbar_mux_001:src_endofpacket -> onchip_memory_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire         cmd_xbar_mux_001_src_valid;                                                                        // cmd_xbar_mux_001:src_valid -> onchip_memory_s1_translator_avalon_universal_slave_0_agent:cp_valid
	wire         cmd_xbar_mux_001_src_startofpacket;                                                                // cmd_xbar_mux_001:src_startofpacket -> onchip_memory_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [75:0] cmd_xbar_mux_001_src_data;                                                                         // cmd_xbar_mux_001:src_data -> onchip_memory_s1_translator_avalon_universal_slave_0_agent:cp_data
	wire  [13:0] cmd_xbar_mux_001_src_channel;                                                                      // cmd_xbar_mux_001:src_channel -> onchip_memory_s1_translator_avalon_universal_slave_0_agent:cp_channel
	wire         cmd_xbar_mux_001_src_ready;                                                                        // onchip_memory_s1_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_mux_001:src_ready
	wire         id_router_001_src_endofpacket;                                                                     // id_router_001:src_endofpacket -> rsp_xbar_demux_001:sink_endofpacket
	wire         id_router_001_src_valid;                                                                           // id_router_001:src_valid -> rsp_xbar_demux_001:sink_valid
	wire         id_router_001_src_startofpacket;                                                                   // id_router_001:src_startofpacket -> rsp_xbar_demux_001:sink_startofpacket
	wire  [75:0] id_router_001_src_data;                                                                            // id_router_001:src_data -> rsp_xbar_demux_001:sink_data
	wire  [13:0] id_router_001_src_channel;                                                                         // id_router_001:src_channel -> rsp_xbar_demux_001:sink_channel
	wire         id_router_001_src_ready;                                                                           // rsp_xbar_demux_001:sink_ready -> id_router_001:src_ready
	wire         cmd_xbar_demux_001_src2_ready;                                                                     // jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_001:src2_ready
	wire         id_router_002_src_endofpacket;                                                                     // id_router_002:src_endofpacket -> rsp_xbar_demux_002:sink_endofpacket
	wire         id_router_002_src_valid;                                                                           // id_router_002:src_valid -> rsp_xbar_demux_002:sink_valid
	wire         id_router_002_src_startofpacket;                                                                   // id_router_002:src_startofpacket -> rsp_xbar_demux_002:sink_startofpacket
	wire  [75:0] id_router_002_src_data;                                                                            // id_router_002:src_data -> rsp_xbar_demux_002:sink_data
	wire  [13:0] id_router_002_src_channel;                                                                         // id_router_002:src_channel -> rsp_xbar_demux_002:sink_channel
	wire         id_router_002_src_ready;                                                                           // rsp_xbar_demux_002:sink_ready -> id_router_002:src_ready
	wire         cmd_xbar_demux_001_src3_ready;                                                                     // sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_001:src3_ready
	wire         id_router_003_src_endofpacket;                                                                     // id_router_003:src_endofpacket -> rsp_xbar_demux_003:sink_endofpacket
	wire         id_router_003_src_valid;                                                                           // id_router_003:src_valid -> rsp_xbar_demux_003:sink_valid
	wire         id_router_003_src_startofpacket;                                                                   // id_router_003:src_startofpacket -> rsp_xbar_demux_003:sink_startofpacket
	wire  [75:0] id_router_003_src_data;                                                                            // id_router_003:src_data -> rsp_xbar_demux_003:sink_data
	wire  [13:0] id_router_003_src_channel;                                                                         // id_router_003:src_channel -> rsp_xbar_demux_003:sink_channel
	wire         id_router_003_src_ready;                                                                           // rsp_xbar_demux_003:sink_ready -> id_router_003:src_ready
	wire         cmd_xbar_demux_001_src4_ready;                                                                     // pio_LEDG_s1_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_001:src4_ready
	wire         id_router_004_src_endofpacket;                                                                     // id_router_004:src_endofpacket -> rsp_xbar_demux_004:sink_endofpacket
	wire         id_router_004_src_valid;                                                                           // id_router_004:src_valid -> rsp_xbar_demux_004:sink_valid
	wire         id_router_004_src_startofpacket;                                                                   // id_router_004:src_startofpacket -> rsp_xbar_demux_004:sink_startofpacket
	wire  [75:0] id_router_004_src_data;                                                                            // id_router_004:src_data -> rsp_xbar_demux_004:sink_data
	wire  [13:0] id_router_004_src_channel;                                                                         // id_router_004:src_channel -> rsp_xbar_demux_004:sink_channel
	wire         id_router_004_src_ready;                                                                           // rsp_xbar_demux_004:sink_ready -> id_router_004:src_ready
	wire         cmd_xbar_demux_001_src5_ready;                                                                     // pio_LEDR_s1_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_001:src5_ready
	wire         id_router_005_src_endofpacket;                                                                     // id_router_005:src_endofpacket -> rsp_xbar_demux_005:sink_endofpacket
	wire         id_router_005_src_valid;                                                                           // id_router_005:src_valid -> rsp_xbar_demux_005:sink_valid
	wire         id_router_005_src_startofpacket;                                                                   // id_router_005:src_startofpacket -> rsp_xbar_demux_005:sink_startofpacket
	wire  [75:0] id_router_005_src_data;                                                                            // id_router_005:src_data -> rsp_xbar_demux_005:sink_data
	wire  [13:0] id_router_005_src_channel;                                                                         // id_router_005:src_channel -> rsp_xbar_demux_005:sink_channel
	wire         id_router_005_src_ready;                                                                           // rsp_xbar_demux_005:sink_ready -> id_router_005:src_ready
	wire         cmd_xbar_demux_001_src6_ready;                                                                     // pio_SW_s1_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_001:src6_ready
	wire         id_router_006_src_endofpacket;                                                                     // id_router_006:src_endofpacket -> rsp_xbar_demux_006:sink_endofpacket
	wire         id_router_006_src_valid;                                                                           // id_router_006:src_valid -> rsp_xbar_demux_006:sink_valid
	wire         id_router_006_src_startofpacket;                                                                   // id_router_006:src_startofpacket -> rsp_xbar_demux_006:sink_startofpacket
	wire  [75:0] id_router_006_src_data;                                                                            // id_router_006:src_data -> rsp_xbar_demux_006:sink_data
	wire  [13:0] id_router_006_src_channel;                                                                         // id_router_006:src_channel -> rsp_xbar_demux_006:sink_channel
	wire         id_router_006_src_ready;                                                                           // rsp_xbar_demux_006:sink_ready -> id_router_006:src_ready
	wire         cmd_xbar_demux_001_src7_ready;                                                                     // pio_Button_s1_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_001:src7_ready
	wire         id_router_007_src_endofpacket;                                                                     // id_router_007:src_endofpacket -> rsp_xbar_demux_007:sink_endofpacket
	wire         id_router_007_src_valid;                                                                           // id_router_007:src_valid -> rsp_xbar_demux_007:sink_valid
	wire         id_router_007_src_startofpacket;                                                                   // id_router_007:src_startofpacket -> rsp_xbar_demux_007:sink_startofpacket
	wire  [75:0] id_router_007_src_data;                                                                            // id_router_007:src_data -> rsp_xbar_demux_007:sink_data
	wire  [13:0] id_router_007_src_channel;                                                                         // id_router_007:src_channel -> rsp_xbar_demux_007:sink_channel
	wire         id_router_007_src_ready;                                                                           // rsp_xbar_demux_007:sink_ready -> id_router_007:src_ready
	wire         cmd_xbar_demux_001_src8_ready;                                                                     // lcd_control_slave_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_001:src8_ready
	wire         id_router_008_src_endofpacket;                                                                     // id_router_008:src_endofpacket -> rsp_xbar_demux_008:sink_endofpacket
	wire         id_router_008_src_valid;                                                                           // id_router_008:src_valid -> rsp_xbar_demux_008:sink_valid
	wire         id_router_008_src_startofpacket;                                                                   // id_router_008:src_startofpacket -> rsp_xbar_demux_008:sink_startofpacket
	wire  [75:0] id_router_008_src_data;                                                                            // id_router_008:src_data -> rsp_xbar_demux_008:sink_data
	wire  [13:0] id_router_008_src_channel;                                                                         // id_router_008:src_channel -> rsp_xbar_demux_008:sink_channel
	wire         id_router_008_src_ready;                                                                           // rsp_xbar_demux_008:sink_ready -> id_router_008:src_ready
	wire         cmd_xbar_demux_001_src9_ready;                                                                     // uart_s1_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_001:src9_ready
	wire         id_router_009_src_endofpacket;                                                                     // id_router_009:src_endofpacket -> rsp_xbar_demux_009:sink_endofpacket
	wire         id_router_009_src_valid;                                                                           // id_router_009:src_valid -> rsp_xbar_demux_009:sink_valid
	wire         id_router_009_src_startofpacket;                                                                   // id_router_009:src_startofpacket -> rsp_xbar_demux_009:sink_startofpacket
	wire  [75:0] id_router_009_src_data;                                                                            // id_router_009:src_data -> rsp_xbar_demux_009:sink_data
	wire  [13:0] id_router_009_src_channel;                                                                         // id_router_009:src_channel -> rsp_xbar_demux_009:sink_channel
	wire         id_router_009_src_ready;                                                                           // rsp_xbar_demux_009:sink_ready -> id_router_009:src_ready
	wire         cmd_xbar_demux_001_src10_ready;                                                                    // timer_0_s1_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_001:src10_ready
	wire         id_router_010_src_endofpacket;                                                                     // id_router_010:src_endofpacket -> rsp_xbar_demux_010:sink_endofpacket
	wire         id_router_010_src_valid;                                                                           // id_router_010:src_valid -> rsp_xbar_demux_010:sink_valid
	wire         id_router_010_src_startofpacket;                                                                   // id_router_010:src_startofpacket -> rsp_xbar_demux_010:sink_startofpacket
	wire  [75:0] id_router_010_src_data;                                                                            // id_router_010:src_data -> rsp_xbar_demux_010:sink_data
	wire  [13:0] id_router_010_src_channel;                                                                         // id_router_010:src_channel -> rsp_xbar_demux_010:sink_channel
	wire         id_router_010_src_ready;                                                                           // rsp_xbar_demux_010:sink_ready -> id_router_010:src_ready
	wire         cmd_xbar_demux_001_src11_ready;                                                                    // pio_Data_s1_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_001:src11_ready
	wire         id_router_011_src_endofpacket;                                                                     // id_router_011:src_endofpacket -> rsp_xbar_demux_011:sink_endofpacket
	wire         id_router_011_src_valid;                                                                           // id_router_011:src_valid -> rsp_xbar_demux_011:sink_valid
	wire         id_router_011_src_startofpacket;                                                                   // id_router_011:src_startofpacket -> rsp_xbar_demux_011:sink_startofpacket
	wire  [75:0] id_router_011_src_data;                                                                            // id_router_011:src_data -> rsp_xbar_demux_011:sink_data
	wire  [13:0] id_router_011_src_channel;                                                                         // id_router_011:src_channel -> rsp_xbar_demux_011:sink_channel
	wire         id_router_011_src_ready;                                                                           // rsp_xbar_demux_011:sink_ready -> id_router_011:src_ready
	wire         cmd_xbar_demux_001_src12_ready;                                                                    // pio_RdyData_s1_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_001:src12_ready
	wire         id_router_012_src_endofpacket;                                                                     // id_router_012:src_endofpacket -> rsp_xbar_demux_012:sink_endofpacket
	wire         id_router_012_src_valid;                                                                           // id_router_012:src_valid -> rsp_xbar_demux_012:sink_valid
	wire         id_router_012_src_startofpacket;                                                                   // id_router_012:src_startofpacket -> rsp_xbar_demux_012:sink_startofpacket
	wire  [75:0] id_router_012_src_data;                                                                            // id_router_012:src_data -> rsp_xbar_demux_012:sink_data
	wire  [13:0] id_router_012_src_channel;                                                                         // id_router_012:src_channel -> rsp_xbar_demux_012:sink_channel
	wire         id_router_012_src_ready;                                                                           // rsp_xbar_demux_012:sink_ready -> id_router_012:src_ready
	wire         cmd_xbar_demux_001_src13_ready;                                                                    // pio_DataRead_s1_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_001:src13_ready
	wire         id_router_013_src_endofpacket;                                                                     // id_router_013:src_endofpacket -> rsp_xbar_demux_013:sink_endofpacket
	wire         id_router_013_src_valid;                                                                           // id_router_013:src_valid -> rsp_xbar_demux_013:sink_valid
	wire         id_router_013_src_startofpacket;                                                                   // id_router_013:src_startofpacket -> rsp_xbar_demux_013:sink_startofpacket
	wire  [75:0] id_router_013_src_data;                                                                            // id_router_013:src_data -> rsp_xbar_demux_013:sink_data
	wire  [13:0] id_router_013_src_channel;                                                                         // id_router_013:src_channel -> rsp_xbar_demux_013:sink_channel
	wire         id_router_013_src_ready;                                                                           // rsp_xbar_demux_013:sink_ready -> id_router_013:src_ready
	wire  [13:0] limiter_cmd_valid_data;                                                                            // limiter:cmd_src_valid -> cmd_xbar_demux:sink_valid
	wire  [13:0] limiter_001_cmd_valid_data;                                                                        // limiter_001:cmd_src_valid -> cmd_xbar_demux_001:sink_valid
	wire         irq_mapper_receiver0_irq;                                                                          // jtag_uart:av_irq -> irq_mapper:receiver0_irq
	wire         irq_mapper_receiver1_irq;                                                                          // timer_0:irq -> irq_mapper:receiver1_irq
	wire         irq_mapper_receiver2_irq;                                                                          // uart:irq -> irq_mapper:receiver2_irq
	wire         irq_mapper_receiver3_irq;                                                                          // pio_Button:irq -> irq_mapper:receiver3_irq
	wire         irq_mapper_receiver4_irq;                                                                          // pio_RdyData:irq -> irq_mapper:receiver4_irq
	wire  [31:0] nios2_qsys_d_irq_irq;                                                                              // irq_mapper:sender_irq -> nios2_qsys:d_irq

	Nios1_nios2_qsys nios2_qsys (
		.clk                                   (clk_clk),                                                                   //                       clk.clk
		.reset_n                               (~rst_controller_reset_out_reset),                                           //                   reset_n.reset_n
		.d_address                             (nios2_qsys_data_master_address),                                            //               data_master.address
		.d_byteenable                          (nios2_qsys_data_master_byteenable),                                         //                          .byteenable
		.d_read                                (nios2_qsys_data_master_read),                                               //                          .read
		.d_readdata                            (nios2_qsys_data_master_readdata),                                           //                          .readdata
		.d_waitrequest                         (nios2_qsys_data_master_waitrequest),                                        //                          .waitrequest
		.d_write                               (nios2_qsys_data_master_write),                                              //                          .write
		.d_writedata                           (nios2_qsys_data_master_writedata),                                          //                          .writedata
		.d_readdatavalid                       (nios2_qsys_data_master_readdatavalid),                                      //                          .readdatavalid
		.jtag_debug_module_debugaccess_to_roms (nios2_qsys_data_master_debugaccess),                                        //                          .debugaccess
		.i_address                             (nios2_qsys_instruction_master_address),                                     //        instruction_master.address
		.i_read                                (nios2_qsys_instruction_master_read),                                        //                          .read
		.i_readdata                            (nios2_qsys_instruction_master_readdata),                                    //                          .readdata
		.i_waitrequest                         (nios2_qsys_instruction_master_waitrequest),                                 //                          .waitrequest
		.i_readdatavalid                       (nios2_qsys_instruction_master_readdatavalid),                               //                          .readdatavalid
		.d_irq                                 (nios2_qsys_d_irq_irq),                                                      //                     d_irq.irq
		.jtag_debug_module_resetrequest        (),                                                                          //   jtag_debug_module_reset.reset
		.jtag_debug_module_address             (nios2_qsys_jtag_debug_module_translator_avalon_anti_slave_0_address),       //         jtag_debug_module.address
		.jtag_debug_module_begintransfer       (nios2_qsys_jtag_debug_module_translator_avalon_anti_slave_0_begintransfer), //                          .begintransfer
		.jtag_debug_module_byteenable          (nios2_qsys_jtag_debug_module_translator_avalon_anti_slave_0_byteenable),    //                          .byteenable
		.jtag_debug_module_debugaccess         (nios2_qsys_jtag_debug_module_translator_avalon_anti_slave_0_debugaccess),   //                          .debugaccess
		.jtag_debug_module_readdata            (nios2_qsys_jtag_debug_module_translator_avalon_anti_slave_0_readdata),      //                          .readdata
		.jtag_debug_module_select              (nios2_qsys_jtag_debug_module_translator_avalon_anti_slave_0_chipselect),    //                          .chipselect
		.jtag_debug_module_write               (nios2_qsys_jtag_debug_module_translator_avalon_anti_slave_0_write),         //                          .write
		.jtag_debug_module_writedata           (nios2_qsys_jtag_debug_module_translator_avalon_anti_slave_0_writedata),     //                          .writedata
		.no_ci_readra                          ()                                                                           // custom_instruction_master.readra
	);

	Nios1_onchip_memory onchip_memory (
		.clk        (clk_clk),                                                    //   clk1.clk
		.address    (onchip_memory_s1_translator_avalon_anti_slave_0_address),    //     s1.address
		.chipselect (onchip_memory_s1_translator_avalon_anti_slave_0_chipselect), //       .chipselect
		.clken      (onchip_memory_s1_translator_avalon_anti_slave_0_clken),      //       .clken
		.readdata   (onchip_memory_s1_translator_avalon_anti_slave_0_readdata),   //       .readdata
		.write      (onchip_memory_s1_translator_avalon_anti_slave_0_write),      //       .write
		.writedata  (onchip_memory_s1_translator_avalon_anti_slave_0_writedata),  //       .writedata
		.byteenable (onchip_memory_s1_translator_avalon_anti_slave_0_byteenable), //       .byteenable
		.reset      (rst_controller_reset_out_reset)                              // reset1.reset
	);

	Nios1_jtag_uart jtag_uart (
		.clk            (clk_clk),                                                                //               clk.clk
		.rst_n          (~rst_controller_reset_out_reset),                                        //             reset.reset_n
		.av_chipselect  (jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_chipselect),  // avalon_jtag_slave.chipselect
		.av_address     (jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_address),     //                  .address
		.av_read_n      (~jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_read),       //                  .read_n
		.av_readdata    (jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_readdata),    //                  .readdata
		.av_write_n     (~jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_write),      //                  .write_n
		.av_writedata   (jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_writedata),   //                  .writedata
		.av_waitrequest (jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_waitrequest), //                  .waitrequest
		.dataavailable  (),                                                                       //                  .dataavailable
		.readyfordata   (),                                                                       //                  .readyfordata
		.av_irq         (irq_mapper_receiver0_irq)                                                //               irq.irq
	);

	Nios1_sysid_qsys sysid_qsys (
		.clock    (clk_clk),                                                          //           clk.clk
		.reset_n  (~rst_controller_reset_out_reset),                                  //         reset.reset_n
		.readdata (sysid_qsys_control_slave_translator_avalon_anti_slave_0_readdata), // control_slave.readdata
		.address  (sysid_qsys_control_slave_translator_avalon_anti_slave_0_address)   //              .address
	);

	Nios1_pio_LEDG pio_ledg (
		.clk        (clk_clk),                                               //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),                       //               reset.reset_n
		.address    (pio_ledg_s1_translator_avalon_anti_slave_0_address),    //                  s1.address
		.write_n    (~pio_ledg_s1_translator_avalon_anti_slave_0_write),     //                    .write_n
		.writedata  (pio_ledg_s1_translator_avalon_anti_slave_0_writedata),  //                    .writedata
		.chipselect (pio_ledg_s1_translator_avalon_anti_slave_0_chipselect), //                    .chipselect
		.readdata   (pio_ledg_s1_translator_avalon_anti_slave_0_readdata),   //                    .readdata
		.out_port   (pio_ledg_export)                                        // external_connection.export
	);

	Nios1_pio_LEDR pio_ledr (
		.clk        (clk_clk),                                               //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),                       //               reset.reset_n
		.address    (pio_ledr_s1_translator_avalon_anti_slave_0_address),    //                  s1.address
		.write_n    (~pio_ledr_s1_translator_avalon_anti_slave_0_write),     //                    .write_n
		.writedata  (pio_ledr_s1_translator_avalon_anti_slave_0_writedata),  //                    .writedata
		.chipselect (pio_ledr_s1_translator_avalon_anti_slave_0_chipselect), //                    .chipselect
		.readdata   (pio_ledr_s1_translator_avalon_anti_slave_0_readdata),   //                    .readdata
		.out_port   (pio_ledr_export)                                        // external_connection.export
	);

	Nios1_pio_SW pio_sw (
		.clk      (clk_clk),                                           //                 clk.clk
		.reset_n  (~rst_controller_reset_out_reset),                   //               reset.reset_n
		.address  (pio_sw_s1_translator_avalon_anti_slave_0_address),  //                  s1.address
		.readdata (pio_sw_s1_translator_avalon_anti_slave_0_readdata), //                    .readdata
		.in_port  (pio_sw_export)                                      // external_connection.export
	);

	Nios1_pio_Button pio_button (
		.clk        (clk_clk),                                                 //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),                         //               reset.reset_n
		.address    (pio_button_s1_translator_avalon_anti_slave_0_address),    //                  s1.address
		.write_n    (~pio_button_s1_translator_avalon_anti_slave_0_write),     //                    .write_n
		.writedata  (pio_button_s1_translator_avalon_anti_slave_0_writedata),  //                    .writedata
		.chipselect (pio_button_s1_translator_avalon_anti_slave_0_chipselect), //                    .chipselect
		.readdata   (pio_button_s1_translator_avalon_anti_slave_0_readdata),   //                    .readdata
		.in_port    (pio_button_export),                                       // external_connection.export
		.irq        (irq_mapper_receiver3_irq)                                 //                 irq.irq
	);

	Nios1_lcd lcd (
		.clk           (clk_clk),                                                        //           clk.clk
		.reset_n       (~rst_controller_reset_out_reset),                                //         reset.reset_n
		.address       (lcd_control_slave_translator_avalon_anti_slave_0_address),       // control_slave.address
		.begintransfer (lcd_control_slave_translator_avalon_anti_slave_0_begintransfer), //              .begintransfer
		.read          (lcd_control_slave_translator_avalon_anti_slave_0_read),          //              .read
		.readdata      (lcd_control_slave_translator_avalon_anti_slave_0_readdata),      //              .readdata
		.write         (lcd_control_slave_translator_avalon_anti_slave_0_write),         //              .write
		.writedata     (lcd_control_slave_translator_avalon_anti_slave_0_writedata),     //              .writedata
		.LCD_data      (lcd_external_data),                                              //      external.export
		.LCD_E         (lcd_external_E),                                                 //              .export
		.LCD_RS        (lcd_external_RS),                                                //              .export
		.LCD_RW        (lcd_external_RW)                                                 //              .export
	);

	Nios1_uart uart (
		.clk           (clk_clk),                                              //                 clk.clk
		.reset_n       (~rst_controller_reset_out_reset),                      //               reset.reset_n
		.address       (uart_s1_translator_avalon_anti_slave_0_address),       //                  s1.address
		.begintransfer (uart_s1_translator_avalon_anti_slave_0_begintransfer), //                    .begintransfer
		.chipselect    (uart_s1_translator_avalon_anti_slave_0_chipselect),    //                    .chipselect
		.read_n        (~uart_s1_translator_avalon_anti_slave_0_read),         //                    .read_n
		.write_n       (~uart_s1_translator_avalon_anti_slave_0_write),        //                    .write_n
		.writedata     (uart_s1_translator_avalon_anti_slave_0_writedata),     //                    .writedata
		.readdata      (uart_s1_translator_avalon_anti_slave_0_readdata),      //                    .readdata
		.dataavailable (),                                                     //                    .dataavailable
		.readyfordata  (),                                                     //                    .readyfordata
		.rxd           (uart_external_rxd),                                    // external_connection.export
		.txd           (uart_external_txd),                                    //                    .export
		.irq           (irq_mapper_receiver2_irq)                              //                 irq.irq
	);

	Nios1_timer_0 timer_0 (
		.clk        (clk_clk),                                              //   clk.clk
		.reset_n    (~rst_controller_reset_out_reset),                      // reset.reset_n
		.address    (timer_0_s1_translator_avalon_anti_slave_0_address),    //    s1.address
		.writedata  (timer_0_s1_translator_avalon_anti_slave_0_writedata),  //      .writedata
		.readdata   (timer_0_s1_translator_avalon_anti_slave_0_readdata),   //      .readdata
		.chipselect (timer_0_s1_translator_avalon_anti_slave_0_chipselect), //      .chipselect
		.write_n    (~timer_0_s1_translator_avalon_anti_slave_0_write),     //      .write_n
		.irq        (irq_mapper_receiver1_irq)                              //   irq.irq
	);

	Nios1_pio_Data pio_data (
		.clk      (clk_clk),                                             //                 clk.clk
		.reset_n  (~rst_controller_reset_out_reset),                     //               reset.reset_n
		.address  (pio_data_s1_translator_avalon_anti_slave_0_address),  //                  s1.address
		.readdata (pio_data_s1_translator_avalon_anti_slave_0_readdata), //                    .readdata
		.in_port  (pio_data_export)                                      // external_connection.export
	);

	Nios1_pio_RdyData pio_rdydata (
		.clk        (clk_clk),                                                  //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),                          //               reset.reset_n
		.address    (pio_rdydata_s1_translator_avalon_anti_slave_0_address),    //                  s1.address
		.write_n    (~pio_rdydata_s1_translator_avalon_anti_slave_0_write),     //                    .write_n
		.writedata  (pio_rdydata_s1_translator_avalon_anti_slave_0_writedata),  //                    .writedata
		.chipselect (pio_rdydata_s1_translator_avalon_anti_slave_0_chipselect), //                    .chipselect
		.readdata   (pio_rdydata_s1_translator_avalon_anti_slave_0_readdata),   //                    .readdata
		.in_port    (pio_rdydata_export),                                       // external_connection.export
		.irq        (irq_mapper_receiver4_irq)                                  //                 irq.irq
	);

	Nios1_pio_DataRead pio_dataread (
		.clk        (clk_clk),                                                   //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),                           //               reset.reset_n
		.address    (pio_dataread_s1_translator_avalon_anti_slave_0_address),    //                  s1.address
		.write_n    (~pio_dataread_s1_translator_avalon_anti_slave_0_write),     //                    .write_n
		.writedata  (pio_dataread_s1_translator_avalon_anti_slave_0_writedata),  //                    .writedata
		.chipselect (pio_dataread_s1_translator_avalon_anti_slave_0_chipselect), //                    .chipselect
		.readdata   (pio_dataread_s1_translator_avalon_anti_slave_0_readdata),   //                    .readdata
		.out_port   (pio_dataread_export)                                        // external_connection.export
	);

	altera_merlin_master_translator #(
		.AV_ADDRESS_W                (19),
		.AV_DATA_W                   (32),
		.AV_BURSTCOUNT_W             (1),
		.AV_BYTEENABLE_W             (4),
		.UAV_ADDRESS_W               (19),
		.UAV_BURSTCOUNT_W            (3),
		.USE_READ                    (1),
		.USE_WRITE                   (0),
		.USE_BEGINBURSTTRANSFER      (0),
		.USE_BEGINTRANSFER           (0),
		.USE_CHIPSELECT              (0),
		.USE_BURSTCOUNT              (0),
		.USE_READDATAVALID           (1),
		.USE_WAITREQUEST             (1),
		.AV_SYMBOLS_PER_WORD         (4),
		.AV_ADDRESS_SYMBOLS          (1),
		.AV_BURSTCOUNT_SYMBOLS       (0),
		.AV_CONSTANT_BURST_BEHAVIOR  (0),
		.UAV_CONSTANT_BURST_BEHAVIOR (0),
		.AV_LINEWRAPBURSTS           (1),
		.AV_REGISTERINCOMINGSIGNALS  (0)
	) nios2_qsys_instruction_master_translator (
		.clk                   (clk_clk),                                                                          //                       clk.clk
		.reset                 (rst_controller_reset_out_reset),                                                   //                     reset.reset
		.uav_address           (nios2_qsys_instruction_master_translator_avalon_universal_master_0_address),       // avalon_universal_master_0.address
		.uav_burstcount        (nios2_qsys_instruction_master_translator_avalon_universal_master_0_burstcount),    //                          .burstcount
		.uav_read              (nios2_qsys_instruction_master_translator_avalon_universal_master_0_read),          //                          .read
		.uav_write             (nios2_qsys_instruction_master_translator_avalon_universal_master_0_write),         //                          .write
		.uav_waitrequest       (nios2_qsys_instruction_master_translator_avalon_universal_master_0_waitrequest),   //                          .waitrequest
		.uav_readdatavalid     (nios2_qsys_instruction_master_translator_avalon_universal_master_0_readdatavalid), //                          .readdatavalid
		.uav_byteenable        (nios2_qsys_instruction_master_translator_avalon_universal_master_0_byteenable),    //                          .byteenable
		.uav_readdata          (nios2_qsys_instruction_master_translator_avalon_universal_master_0_readdata),      //                          .readdata
		.uav_writedata         (nios2_qsys_instruction_master_translator_avalon_universal_master_0_writedata),     //                          .writedata
		.uav_lock              (nios2_qsys_instruction_master_translator_avalon_universal_master_0_lock),          //                          .lock
		.uav_debugaccess       (nios2_qsys_instruction_master_translator_avalon_universal_master_0_debugaccess),   //                          .debugaccess
		.av_address            (nios2_qsys_instruction_master_address),                                            //      avalon_anti_master_0.address
		.av_waitrequest        (nios2_qsys_instruction_master_waitrequest),                                        //                          .waitrequest
		.av_read               (nios2_qsys_instruction_master_read),                                               //                          .read
		.av_readdata           (nios2_qsys_instruction_master_readdata),                                           //                          .readdata
		.av_readdatavalid      (nios2_qsys_instruction_master_readdatavalid),                                      //                          .readdatavalid
		.av_burstcount         (1'b1),                                                                             //               (terminated)
		.av_byteenable         (4'b1111),                                                                          //               (terminated)
		.av_beginbursttransfer (1'b0),                                                                             //               (terminated)
		.av_begintransfer      (1'b0),                                                                             //               (terminated)
		.av_chipselect         (1'b0),                                                                             //               (terminated)
		.av_write              (1'b0),                                                                             //               (terminated)
		.av_writedata          (32'b00000000000000000000000000000000),                                             //               (terminated)
		.av_lock               (1'b0),                                                                             //               (terminated)
		.av_debugaccess        (1'b0),                                                                             //               (terminated)
		.uav_clken             (),                                                                                 //               (terminated)
		.av_clken              (1'b1)                                                                              //               (terminated)
	);

	altera_merlin_master_translator #(
		.AV_ADDRESS_W                (19),
		.AV_DATA_W                   (32),
		.AV_BURSTCOUNT_W             (1),
		.AV_BYTEENABLE_W             (4),
		.UAV_ADDRESS_W               (19),
		.UAV_BURSTCOUNT_W            (3),
		.USE_READ                    (1),
		.USE_WRITE                   (1),
		.USE_BEGINBURSTTRANSFER      (0),
		.USE_BEGINTRANSFER           (0),
		.USE_CHIPSELECT              (0),
		.USE_BURSTCOUNT              (0),
		.USE_READDATAVALID           (1),
		.USE_WAITREQUEST             (1),
		.AV_SYMBOLS_PER_WORD         (4),
		.AV_ADDRESS_SYMBOLS          (1),
		.AV_BURSTCOUNT_SYMBOLS       (0),
		.AV_CONSTANT_BURST_BEHAVIOR  (0),
		.UAV_CONSTANT_BURST_BEHAVIOR (0),
		.AV_LINEWRAPBURSTS           (0),
		.AV_REGISTERINCOMINGSIGNALS  (0)
	) nios2_qsys_data_master_translator (
		.clk                   (clk_clk),                                                                   //                       clk.clk
		.reset                 (rst_controller_reset_out_reset),                                            //                     reset.reset
		.uav_address           (nios2_qsys_data_master_translator_avalon_universal_master_0_address),       // avalon_universal_master_0.address
		.uav_burstcount        (nios2_qsys_data_master_translator_avalon_universal_master_0_burstcount),    //                          .burstcount
		.uav_read              (nios2_qsys_data_master_translator_avalon_universal_master_0_read),          //                          .read
		.uav_write             (nios2_qsys_data_master_translator_avalon_universal_master_0_write),         //                          .write
		.uav_waitrequest       (nios2_qsys_data_master_translator_avalon_universal_master_0_waitrequest),   //                          .waitrequest
		.uav_readdatavalid     (nios2_qsys_data_master_translator_avalon_universal_master_0_readdatavalid), //                          .readdatavalid
		.uav_byteenable        (nios2_qsys_data_master_translator_avalon_universal_master_0_byteenable),    //                          .byteenable
		.uav_readdata          (nios2_qsys_data_master_translator_avalon_universal_master_0_readdata),      //                          .readdata
		.uav_writedata         (nios2_qsys_data_master_translator_avalon_universal_master_0_writedata),     //                          .writedata
		.uav_lock              (nios2_qsys_data_master_translator_avalon_universal_master_0_lock),          //                          .lock
		.uav_debugaccess       (nios2_qsys_data_master_translator_avalon_universal_master_0_debugaccess),   //                          .debugaccess
		.av_address            (nios2_qsys_data_master_address),                                            //      avalon_anti_master_0.address
		.av_waitrequest        (nios2_qsys_data_master_waitrequest),                                        //                          .waitrequest
		.av_byteenable         (nios2_qsys_data_master_byteenable),                                         //                          .byteenable
		.av_read               (nios2_qsys_data_master_read),                                               //                          .read
		.av_readdata           (nios2_qsys_data_master_readdata),                                           //                          .readdata
		.av_readdatavalid      (nios2_qsys_data_master_readdatavalid),                                      //                          .readdatavalid
		.av_write              (nios2_qsys_data_master_write),                                              //                          .write
		.av_writedata          (nios2_qsys_data_master_writedata),                                          //                          .writedata
		.av_debugaccess        (nios2_qsys_data_master_debugaccess),                                        //                          .debugaccess
		.av_burstcount         (1'b1),                                                                      //               (terminated)
		.av_beginbursttransfer (1'b0),                                                                      //               (terminated)
		.av_begintransfer      (1'b0),                                                                      //               (terminated)
		.av_chipselect         (1'b0),                                                                      //               (terminated)
		.av_lock               (1'b0),                                                                      //               (terminated)
		.uav_clken             (),                                                                          //               (terminated)
		.av_clken              (1'b1)                                                                       //               (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (9),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (4),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (19),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) nios2_qsys_jtag_debug_module_translator (
		.clk                   (clk_clk),                                                                                 //                      clk.clk
		.reset                 (rst_controller_reset_out_reset),                                                          //                    reset.reset
		.uav_address           (nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount        (nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read              (nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write             (nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest       (nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid     (nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable        (nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata          (nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata         (nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock              (nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess       (nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address            (nios2_qsys_jtag_debug_module_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write              (nios2_qsys_jtag_debug_module_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_readdata           (nios2_qsys_jtag_debug_module_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata          (nios2_qsys_jtag_debug_module_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_begintransfer      (nios2_qsys_jtag_debug_module_translator_avalon_anti_slave_0_begintransfer),               //                         .begintransfer
		.av_byteenable         (nios2_qsys_jtag_debug_module_translator_avalon_anti_slave_0_byteenable),                  //                         .byteenable
		.av_chipselect         (nios2_qsys_jtag_debug_module_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_debugaccess        (nios2_qsys_jtag_debug_module_translator_avalon_anti_slave_0_debugaccess),                 //                         .debugaccess
		.av_read               (),                                                                                        //              (terminated)
		.av_beginbursttransfer (),                                                                                        //              (terminated)
		.av_burstcount         (),                                                                                        //              (terminated)
		.av_readdatavalid      (1'b0),                                                                                    //              (terminated)
		.av_waitrequest        (1'b0),                                                                                    //              (terminated)
		.av_writebyteenable    (),                                                                                        //              (terminated)
		.av_lock               (),                                                                                        //              (terminated)
		.av_clken              (),                                                                                        //              (terminated)
		.uav_clken             (1'b0),                                                                                    //              (terminated)
		.av_outputenable       ()                                                                                         //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (15),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (4),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (19),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (1),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (0),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) onchip_memory_s1_translator (
		.clk                   (clk_clk),                                                                     //                      clk.clk
		.reset                 (rst_controller_reset_out_reset),                                              //                    reset.reset
		.uav_address           (onchip_memory_s1_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount        (onchip_memory_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read              (onchip_memory_s1_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write             (onchip_memory_s1_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest       (onchip_memory_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid     (onchip_memory_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable        (onchip_memory_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata          (onchip_memory_s1_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata         (onchip_memory_s1_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock              (onchip_memory_s1_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess       (onchip_memory_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address            (onchip_memory_s1_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write              (onchip_memory_s1_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_readdata           (onchip_memory_s1_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata          (onchip_memory_s1_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_byteenable         (onchip_memory_s1_translator_avalon_anti_slave_0_byteenable),                  //                         .byteenable
		.av_chipselect         (onchip_memory_s1_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_clken              (onchip_memory_s1_translator_avalon_anti_slave_0_clken),                       //                         .clken
		.av_read               (),                                                                            //              (terminated)
		.av_begintransfer      (),                                                                            //              (terminated)
		.av_beginbursttransfer (),                                                                            //              (terminated)
		.av_burstcount         (),                                                                            //              (terminated)
		.av_readdatavalid      (1'b0),                                                                        //              (terminated)
		.av_waitrequest        (1'b0),                                                                        //              (terminated)
		.av_writebyteenable    (),                                                                            //              (terminated)
		.av_lock               (),                                                                            //              (terminated)
		.uav_clken             (1'b0),                                                                        //              (terminated)
		.av_debugaccess        (),                                                                            //              (terminated)
		.av_outputenable       ()                                                                             //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (1),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (1),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (19),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (1),
		.USE_UAV_CLKEN                  (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) jtag_uart_avalon_jtag_slave_translator (
		.clk                   (clk_clk),                                                                                //                      clk.clk
		.reset                 (rst_controller_reset_out_reset),                                                         //                    reset.reset
		.uav_address           (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount        (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read              (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write             (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest       (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid     (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable        (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata          (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata         (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock              (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess       (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address            (jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write              (jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_read               (jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_read),                        //                         .read
		.av_readdata           (jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata          (jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_waitrequest        (jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_waitrequest),                 //                         .waitrequest
		.av_chipselect         (jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_begintransfer      (),                                                                                       //              (terminated)
		.av_beginbursttransfer (),                                                                                       //              (terminated)
		.av_burstcount         (),                                                                                       //              (terminated)
		.av_byteenable         (),                                                                                       //              (terminated)
		.av_readdatavalid      (1'b0),                                                                                   //              (terminated)
		.av_writebyteenable    (),                                                                                       //              (terminated)
		.av_lock               (),                                                                                       //              (terminated)
		.av_clken              (),                                                                                       //              (terminated)
		.uav_clken             (1'b0),                                                                                   //              (terminated)
		.av_debugaccess        (),                                                                                       //              (terminated)
		.av_outputenable       ()                                                                                        //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (1),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (4),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (19),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) sysid_qsys_control_slave_translator (
		.clk                   (clk_clk),                                                                             //                      clk.clk
		.reset                 (rst_controller_reset_out_reset),                                                      //                    reset.reset
		.uav_address           (sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount        (sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read              (sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write             (sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest       (sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid     (sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable        (sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata          (sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata         (sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock              (sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess       (sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address            (sysid_qsys_control_slave_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_readdata           (sysid_qsys_control_slave_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_write              (),                                                                                    //              (terminated)
		.av_read               (),                                                                                    //              (terminated)
		.av_writedata          (),                                                                                    //              (terminated)
		.av_begintransfer      (),                                                                                    //              (terminated)
		.av_beginbursttransfer (),                                                                                    //              (terminated)
		.av_burstcount         (),                                                                                    //              (terminated)
		.av_byteenable         (),                                                                                    //              (terminated)
		.av_readdatavalid      (1'b0),                                                                                //              (terminated)
		.av_waitrequest        (1'b0),                                                                                //              (terminated)
		.av_writebyteenable    (),                                                                                    //              (terminated)
		.av_lock               (),                                                                                    //              (terminated)
		.av_chipselect         (),                                                                                    //              (terminated)
		.av_clken              (),                                                                                    //              (terminated)
		.uav_clken             (1'b0),                                                                                //              (terminated)
		.av_debugaccess        (),                                                                                    //              (terminated)
		.av_outputenable       ()                                                                                     //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (3),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (1),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (19),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) pio_ledg_s1_translator (
		.clk                   (clk_clk),                                                                //                      clk.clk
		.reset                 (rst_controller_reset_out_reset),                                         //                    reset.reset
		.uav_address           (pio_ledg_s1_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount        (pio_ledg_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read              (pio_ledg_s1_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write             (pio_ledg_s1_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest       (pio_ledg_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid     (pio_ledg_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable        (pio_ledg_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata          (pio_ledg_s1_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata         (pio_ledg_s1_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock              (pio_ledg_s1_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess       (pio_ledg_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address            (pio_ledg_s1_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write              (pio_ledg_s1_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_readdata           (pio_ledg_s1_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata          (pio_ledg_s1_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_chipselect         (pio_ledg_s1_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_read               (),                                                                       //              (terminated)
		.av_begintransfer      (),                                                                       //              (terminated)
		.av_beginbursttransfer (),                                                                       //              (terminated)
		.av_burstcount         (),                                                                       //              (terminated)
		.av_byteenable         (),                                                                       //              (terminated)
		.av_readdatavalid      (1'b0),                                                                   //              (terminated)
		.av_waitrequest        (1'b0),                                                                   //              (terminated)
		.av_writebyteenable    (),                                                                       //              (terminated)
		.av_lock               (),                                                                       //              (terminated)
		.av_clken              (),                                                                       //              (terminated)
		.uav_clken             (1'b0),                                                                   //              (terminated)
		.av_debugaccess        (),                                                                       //              (terminated)
		.av_outputenable       ()                                                                        //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (3),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (1),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (19),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) pio_ledr_s1_translator (
		.clk                   (clk_clk),                                                                //                      clk.clk
		.reset                 (rst_controller_reset_out_reset),                                         //                    reset.reset
		.uav_address           (pio_ledr_s1_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount        (pio_ledr_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read              (pio_ledr_s1_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write             (pio_ledr_s1_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest       (pio_ledr_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid     (pio_ledr_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable        (pio_ledr_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata          (pio_ledr_s1_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata         (pio_ledr_s1_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock              (pio_ledr_s1_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess       (pio_ledr_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address            (pio_ledr_s1_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write              (pio_ledr_s1_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_readdata           (pio_ledr_s1_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata          (pio_ledr_s1_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_chipselect         (pio_ledr_s1_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_read               (),                                                                       //              (terminated)
		.av_begintransfer      (),                                                                       //              (terminated)
		.av_beginbursttransfer (),                                                                       //              (terminated)
		.av_burstcount         (),                                                                       //              (terminated)
		.av_byteenable         (),                                                                       //              (terminated)
		.av_readdatavalid      (1'b0),                                                                   //              (terminated)
		.av_waitrequest        (1'b0),                                                                   //              (terminated)
		.av_writebyteenable    (),                                                                       //              (terminated)
		.av_lock               (),                                                                       //              (terminated)
		.av_clken              (),                                                                       //              (terminated)
		.uav_clken             (1'b0),                                                                   //              (terminated)
		.av_debugaccess        (),                                                                       //              (terminated)
		.av_outputenable       ()                                                                        //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (2),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (1),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (19),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) pio_sw_s1_translator (
		.clk                   (clk_clk),                                                              //                      clk.clk
		.reset                 (rst_controller_reset_out_reset),                                       //                    reset.reset
		.uav_address           (pio_sw_s1_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount        (pio_sw_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read              (pio_sw_s1_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write             (pio_sw_s1_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest       (pio_sw_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid     (pio_sw_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable        (pio_sw_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata          (pio_sw_s1_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata         (pio_sw_s1_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock              (pio_sw_s1_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess       (pio_sw_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address            (pio_sw_s1_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_readdata           (pio_sw_s1_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_write              (),                                                                     //              (terminated)
		.av_read               (),                                                                     //              (terminated)
		.av_writedata          (),                                                                     //              (terminated)
		.av_begintransfer      (),                                                                     //              (terminated)
		.av_beginbursttransfer (),                                                                     //              (terminated)
		.av_burstcount         (),                                                                     //              (terminated)
		.av_byteenable         (),                                                                     //              (terminated)
		.av_readdatavalid      (1'b0),                                                                 //              (terminated)
		.av_waitrequest        (1'b0),                                                                 //              (terminated)
		.av_writebyteenable    (),                                                                     //              (terminated)
		.av_lock               (),                                                                     //              (terminated)
		.av_chipselect         (),                                                                     //              (terminated)
		.av_clken              (),                                                                     //              (terminated)
		.uav_clken             (1'b0),                                                                 //              (terminated)
		.av_debugaccess        (),                                                                     //              (terminated)
		.av_outputenable       ()                                                                      //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (2),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (1),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (19),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) pio_button_s1_translator (
		.clk                   (clk_clk),                                                                  //                      clk.clk
		.reset                 (rst_controller_reset_out_reset),                                           //                    reset.reset
		.uav_address           (pio_button_s1_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount        (pio_button_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read              (pio_button_s1_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write             (pio_button_s1_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest       (pio_button_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid     (pio_button_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable        (pio_button_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata          (pio_button_s1_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata         (pio_button_s1_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock              (pio_button_s1_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess       (pio_button_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address            (pio_button_s1_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write              (pio_button_s1_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_readdata           (pio_button_s1_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata          (pio_button_s1_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_chipselect         (pio_button_s1_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_read               (),                                                                         //              (terminated)
		.av_begintransfer      (),                                                                         //              (terminated)
		.av_beginbursttransfer (),                                                                         //              (terminated)
		.av_burstcount         (),                                                                         //              (terminated)
		.av_byteenable         (),                                                                         //              (terminated)
		.av_readdatavalid      (1'b0),                                                                     //              (terminated)
		.av_waitrequest        (1'b0),                                                                     //              (terminated)
		.av_writebyteenable    (),                                                                         //              (terminated)
		.av_lock               (),                                                                         //              (terminated)
		.av_clken              (),                                                                         //              (terminated)
		.uav_clken             (1'b0),                                                                     //              (terminated)
		.av_debugaccess        (),                                                                         //              (terminated)
		.av_outputenable       ()                                                                          //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (2),
		.AV_DATA_W                      (8),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (1),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (19),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (13),
		.AV_WRITE_WAIT_CYCLES           (13),
		.AV_SETUP_WAIT_CYCLES           (13),
		.AV_DATA_HOLD_CYCLES            (13)
	) lcd_control_slave_translator (
		.clk                   (clk_clk),                                                                      //                      clk.clk
		.reset                 (rst_controller_reset_out_reset),                                               //                    reset.reset
		.uav_address           (lcd_control_slave_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount        (lcd_control_slave_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read              (lcd_control_slave_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write             (lcd_control_slave_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest       (lcd_control_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid     (lcd_control_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable        (lcd_control_slave_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata          (lcd_control_slave_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata         (lcd_control_slave_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock              (lcd_control_slave_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess       (lcd_control_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address            (lcd_control_slave_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write              (lcd_control_slave_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_read               (lcd_control_slave_translator_avalon_anti_slave_0_read),                        //                         .read
		.av_readdata           (lcd_control_slave_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata          (lcd_control_slave_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_begintransfer      (lcd_control_slave_translator_avalon_anti_slave_0_begintransfer),               //                         .begintransfer
		.av_beginbursttransfer (),                                                                             //              (terminated)
		.av_burstcount         (),                                                                             //              (terminated)
		.av_byteenable         (),                                                                             //              (terminated)
		.av_readdatavalid      (1'b0),                                                                         //              (terminated)
		.av_waitrequest        (1'b0),                                                                         //              (terminated)
		.av_writebyteenable    (),                                                                             //              (terminated)
		.av_lock               (),                                                                             //              (terminated)
		.av_chipselect         (),                                                                             //              (terminated)
		.av_clken              (),                                                                             //              (terminated)
		.uav_clken             (1'b0),                                                                         //              (terminated)
		.av_debugaccess        (),                                                                             //              (terminated)
		.av_outputenable       ()                                                                              //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (3),
		.AV_DATA_W                      (16),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (1),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (19),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (1),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) uart_s1_translator (
		.clk                   (clk_clk),                                                            //                      clk.clk
		.reset                 (rst_controller_reset_out_reset),                                     //                    reset.reset
		.uav_address           (uart_s1_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount        (uart_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read              (uart_s1_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write             (uart_s1_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest       (uart_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid     (uart_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable        (uart_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata          (uart_s1_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata         (uart_s1_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock              (uart_s1_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess       (uart_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address            (uart_s1_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write              (uart_s1_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_read               (uart_s1_translator_avalon_anti_slave_0_read),                        //                         .read
		.av_readdata           (uart_s1_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata          (uart_s1_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_begintransfer      (uart_s1_translator_avalon_anti_slave_0_begintransfer),               //                         .begintransfer
		.av_chipselect         (uart_s1_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_beginbursttransfer (),                                                                   //              (terminated)
		.av_burstcount         (),                                                                   //              (terminated)
		.av_byteenable         (),                                                                   //              (terminated)
		.av_readdatavalid      (1'b0),                                                               //              (terminated)
		.av_waitrequest        (1'b0),                                                               //              (terminated)
		.av_writebyteenable    (),                                                                   //              (terminated)
		.av_lock               (),                                                                   //              (terminated)
		.av_clken              (),                                                                   //              (terminated)
		.uav_clken             (1'b0),                                                               //              (terminated)
		.av_debugaccess        (),                                                                   //              (terminated)
		.av_outputenable       ()                                                                    //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (3),
		.AV_DATA_W                      (16),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (1),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (19),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) timer_0_s1_translator (
		.clk                   (clk_clk),                                                               //                      clk.clk
		.reset                 (rst_controller_reset_out_reset),                                        //                    reset.reset
		.uav_address           (timer_0_s1_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount        (timer_0_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read              (timer_0_s1_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write             (timer_0_s1_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest       (timer_0_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid     (timer_0_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable        (timer_0_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata          (timer_0_s1_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata         (timer_0_s1_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock              (timer_0_s1_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess       (timer_0_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address            (timer_0_s1_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write              (timer_0_s1_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_readdata           (timer_0_s1_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata          (timer_0_s1_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_chipselect         (timer_0_s1_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_read               (),                                                                      //              (terminated)
		.av_begintransfer      (),                                                                      //              (terminated)
		.av_beginbursttransfer (),                                                                      //              (terminated)
		.av_burstcount         (),                                                                      //              (terminated)
		.av_byteenable         (),                                                                      //              (terminated)
		.av_readdatavalid      (1'b0),                                                                  //              (terminated)
		.av_waitrequest        (1'b0),                                                                  //              (terminated)
		.av_writebyteenable    (),                                                                      //              (terminated)
		.av_lock               (),                                                                      //              (terminated)
		.av_clken              (),                                                                      //              (terminated)
		.uav_clken             (1'b0),                                                                  //              (terminated)
		.av_debugaccess        (),                                                                      //              (terminated)
		.av_outputenable       ()                                                                       //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (2),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (1),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (19),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) pio_data_s1_translator (
		.clk                   (clk_clk),                                                                //                      clk.clk
		.reset                 (rst_controller_reset_out_reset),                                         //                    reset.reset
		.uav_address           (pio_data_s1_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount        (pio_data_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read              (pio_data_s1_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write             (pio_data_s1_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest       (pio_data_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid     (pio_data_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable        (pio_data_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata          (pio_data_s1_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata         (pio_data_s1_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock              (pio_data_s1_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess       (pio_data_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address            (pio_data_s1_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_readdata           (pio_data_s1_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_write              (),                                                                       //              (terminated)
		.av_read               (),                                                                       //              (terminated)
		.av_writedata          (),                                                                       //              (terminated)
		.av_begintransfer      (),                                                                       //              (terminated)
		.av_beginbursttransfer (),                                                                       //              (terminated)
		.av_burstcount         (),                                                                       //              (terminated)
		.av_byteenable         (),                                                                       //              (terminated)
		.av_readdatavalid      (1'b0),                                                                   //              (terminated)
		.av_waitrequest        (1'b0),                                                                   //              (terminated)
		.av_writebyteenable    (),                                                                       //              (terminated)
		.av_lock               (),                                                                       //              (terminated)
		.av_chipselect         (),                                                                       //              (terminated)
		.av_clken              (),                                                                       //              (terminated)
		.uav_clken             (1'b0),                                                                   //              (terminated)
		.av_debugaccess        (),                                                                       //              (terminated)
		.av_outputenable       ()                                                                        //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (2),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (1),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (19),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) pio_rdydata_s1_translator (
		.clk                   (clk_clk),                                                                   //                      clk.clk
		.reset                 (rst_controller_reset_out_reset),                                            //                    reset.reset
		.uav_address           (pio_rdydata_s1_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount        (pio_rdydata_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read              (pio_rdydata_s1_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write             (pio_rdydata_s1_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest       (pio_rdydata_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid     (pio_rdydata_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable        (pio_rdydata_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata          (pio_rdydata_s1_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata         (pio_rdydata_s1_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock              (pio_rdydata_s1_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess       (pio_rdydata_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address            (pio_rdydata_s1_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write              (pio_rdydata_s1_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_readdata           (pio_rdydata_s1_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata          (pio_rdydata_s1_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_chipselect         (pio_rdydata_s1_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_read               (),                                                                          //              (terminated)
		.av_begintransfer      (),                                                                          //              (terminated)
		.av_beginbursttransfer (),                                                                          //              (terminated)
		.av_burstcount         (),                                                                          //              (terminated)
		.av_byteenable         (),                                                                          //              (terminated)
		.av_readdatavalid      (1'b0),                                                                      //              (terminated)
		.av_waitrequest        (1'b0),                                                                      //              (terminated)
		.av_writebyteenable    (),                                                                          //              (terminated)
		.av_lock               (),                                                                          //              (terminated)
		.av_clken              (),                                                                          //              (terminated)
		.uav_clken             (1'b0),                                                                      //              (terminated)
		.av_debugaccess        (),                                                                          //              (terminated)
		.av_outputenable       ()                                                                           //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (3),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (1),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (19),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) pio_dataread_s1_translator (
		.clk                   (clk_clk),                                                                    //                      clk.clk
		.reset                 (rst_controller_reset_out_reset),                                             //                    reset.reset
		.uav_address           (pio_dataread_s1_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount        (pio_dataread_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read              (pio_dataread_s1_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write             (pio_dataread_s1_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest       (pio_dataread_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid     (pio_dataread_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable        (pio_dataread_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata          (pio_dataread_s1_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata         (pio_dataread_s1_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock              (pio_dataread_s1_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess       (pio_dataread_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address            (pio_dataread_s1_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write              (pio_dataread_s1_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_readdata           (pio_dataread_s1_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata          (pio_dataread_s1_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_chipselect         (pio_dataread_s1_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_read               (),                                                                           //              (terminated)
		.av_begintransfer      (),                                                                           //              (terminated)
		.av_beginbursttransfer (),                                                                           //              (terminated)
		.av_burstcount         (),                                                                           //              (terminated)
		.av_byteenable         (),                                                                           //              (terminated)
		.av_readdatavalid      (1'b0),                                                                       //              (terminated)
		.av_waitrequest        (1'b0),                                                                       //              (terminated)
		.av_writebyteenable    (),                                                                           //              (terminated)
		.av_lock               (),                                                                           //              (terminated)
		.av_clken              (),                                                                           //              (terminated)
		.uav_clken             (1'b0),                                                                       //              (terminated)
		.av_debugaccess        (),                                                                           //              (terminated)
		.av_outputenable       ()                                                                            //              (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (66),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (54),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (55),
		.PKT_TRANS_POSTED          (56),
		.PKT_TRANS_WRITE           (57),
		.PKT_TRANS_READ            (58),
		.PKT_TRANS_LOCK            (59),
		.PKT_SRC_ID_H              (70),
		.PKT_SRC_ID_L              (67),
		.PKT_DEST_ID_H             (74),
		.PKT_DEST_ID_L             (71),
		.PKT_BURSTWRAP_H           (65),
		.PKT_BURSTWRAP_L           (63),
		.PKT_BYTE_CNT_H            (62),
		.PKT_BYTE_CNT_L            (60),
		.PKT_PROTECTION_H          (75),
		.PKT_PROTECTION_L          (75),
		.ST_CHANNEL_W              (14),
		.ST_DATA_W                 (76),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1)
	) uart_s1_translator_avalon_universal_slave_0_agent (
		.clk                     (clk_clk),                                                                      //             clk.clk
		.reset                   (rst_controller_reset_out_reset),                                               //       clk_reset.reset
		.m0_address              (uart_s1_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (uart_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (uart_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (uart_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (uart_s1_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (uart_s1_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (uart_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (uart_s1_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (uart_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (uart_s1_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (uart_s1_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (uart_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (uart_s1_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (uart_s1_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (uart_s1_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (uart_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_demux_001_src9_ready),                                                //              cp.ready
		.cp_valid                (cmd_xbar_demux_001_src9_valid),                                                //                .valid
		.cp_data                 (cmd_xbar_demux_001_src9_data),                                                 //                .data
		.cp_startofpacket        (cmd_xbar_demux_001_src9_startofpacket),                                        //                .startofpacket
		.cp_endofpacket          (cmd_xbar_demux_001_src9_endofpacket),                                          //                .endofpacket
		.cp_channel              (cmd_xbar_demux_001_src9_channel),                                              //                .channel
		.rf_sink_ready           (uart_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (uart_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (uart_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (uart_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (uart_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (uart_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (uart_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (uart_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (uart_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (uart_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (uart_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (uart_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (uart_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (uart_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (uart_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (uart_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data)         //                .data
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (77),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) uart_s1_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clk_clk),                                                                      //       clk.clk
		.reset             (rst_controller_reset_out_reset),                                               // clk_reset.reset
		.in_data           (uart_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (uart_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (uart_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (uart_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (uart_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (uart_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (uart_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (uart_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (uart_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (uart_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                        // (terminated)
		.csr_read          (1'b0),                                                                         // (terminated)
		.csr_write         (1'b0),                                                                         // (terminated)
		.csr_readdata      (),                                                                             // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                         // (terminated)
		.almost_full_data  (),                                                                             // (terminated)
		.almost_empty_data (),                                                                             // (terminated)
		.in_empty          (1'b0),                                                                         // (terminated)
		.out_empty         (),                                                                             // (terminated)
		.in_error          (1'b0),                                                                         // (terminated)
		.out_error         (),                                                                             // (terminated)
		.in_channel        (1'b0),                                                                         // (terminated)
		.out_channel       ()                                                                              // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (66),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (54),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (55),
		.PKT_TRANS_POSTED          (56),
		.PKT_TRANS_WRITE           (57),
		.PKT_TRANS_READ            (58),
		.PKT_TRANS_LOCK            (59),
		.PKT_SRC_ID_H              (70),
		.PKT_SRC_ID_L              (67),
		.PKT_DEST_ID_H             (74),
		.PKT_DEST_ID_L             (71),
		.PKT_BURSTWRAP_H           (65),
		.PKT_BURSTWRAP_L           (63),
		.PKT_BYTE_CNT_H            (62),
		.PKT_BYTE_CNT_L            (60),
		.PKT_PROTECTION_H          (75),
		.PKT_PROTECTION_L          (75),
		.ST_CHANNEL_W              (14),
		.ST_DATA_W                 (76),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1)
	) pio_dataread_s1_translator_avalon_universal_slave_0_agent (
		.clk                     (clk_clk),                                                                              //             clk.clk
		.reset                   (rst_controller_reset_out_reset),                                                       //       clk_reset.reset
		.m0_address              (pio_dataread_s1_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (pio_dataread_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (pio_dataread_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (pio_dataread_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (pio_dataread_s1_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (pio_dataread_s1_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (pio_dataread_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (pio_dataread_s1_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (pio_dataread_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (pio_dataread_s1_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (pio_dataread_s1_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (pio_dataread_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (pio_dataread_s1_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (pio_dataread_s1_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (pio_dataread_s1_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (pio_dataread_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_demux_001_src13_ready),                                                       //              cp.ready
		.cp_valid                (cmd_xbar_demux_001_src13_valid),                                                       //                .valid
		.cp_data                 (cmd_xbar_demux_001_src13_data),                                                        //                .data
		.cp_startofpacket        (cmd_xbar_demux_001_src13_startofpacket),                                               //                .startofpacket
		.cp_endofpacket          (cmd_xbar_demux_001_src13_endofpacket),                                                 //                .endofpacket
		.cp_channel              (cmd_xbar_demux_001_src13_channel),                                                     //                .channel
		.rf_sink_ready           (pio_dataread_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (pio_dataread_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (pio_dataread_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (pio_dataread_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (pio_dataread_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (pio_dataread_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (pio_dataread_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (pio_dataread_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (pio_dataread_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (pio_dataread_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (pio_dataread_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (pio_dataread_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (pio_dataread_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (pio_dataread_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (pio_dataread_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (pio_dataread_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data)         //                .data
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (77),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) pio_dataread_s1_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clk_clk),                                                                              //       clk.clk
		.reset             (rst_controller_reset_out_reset),                                                       // clk_reset.reset
		.in_data           (pio_dataread_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (pio_dataread_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (pio_dataread_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (pio_dataread_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (pio_dataread_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (pio_dataread_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (pio_dataread_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (pio_dataread_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (pio_dataread_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (pio_dataread_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                // (terminated)
		.csr_read          (1'b0),                                                                                 // (terminated)
		.csr_write         (1'b0),                                                                                 // (terminated)
		.csr_readdata      (),                                                                                     // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                 // (terminated)
		.almost_full_data  (),                                                                                     // (terminated)
		.almost_empty_data (),                                                                                     // (terminated)
		.in_empty          (1'b0),                                                                                 // (terminated)
		.out_empty         (),                                                                                     // (terminated)
		.in_error          (1'b0),                                                                                 // (terminated)
		.out_error         (),                                                                                     // (terminated)
		.in_channel        (1'b0),                                                                                 // (terminated)
		.out_channel       ()                                                                                      // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (66),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (54),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (55),
		.PKT_TRANS_POSTED          (56),
		.PKT_TRANS_WRITE           (57),
		.PKT_TRANS_READ            (58),
		.PKT_TRANS_LOCK            (59),
		.PKT_SRC_ID_H              (70),
		.PKT_SRC_ID_L              (67),
		.PKT_DEST_ID_H             (74),
		.PKT_DEST_ID_L             (71),
		.PKT_BURSTWRAP_H           (65),
		.PKT_BURSTWRAP_L           (63),
		.PKT_BYTE_CNT_H            (62),
		.PKT_BYTE_CNT_L            (60),
		.PKT_PROTECTION_H          (75),
		.PKT_PROTECTION_L          (75),
		.ST_CHANNEL_W              (14),
		.ST_DATA_W                 (76),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1)
	) pio_rdydata_s1_translator_avalon_universal_slave_0_agent (
		.clk                     (clk_clk),                                                                             //             clk.clk
		.reset                   (rst_controller_reset_out_reset),                                                      //       clk_reset.reset
		.m0_address              (pio_rdydata_s1_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (pio_rdydata_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (pio_rdydata_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (pio_rdydata_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (pio_rdydata_s1_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (pio_rdydata_s1_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (pio_rdydata_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (pio_rdydata_s1_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (pio_rdydata_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (pio_rdydata_s1_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (pio_rdydata_s1_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (pio_rdydata_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (pio_rdydata_s1_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (pio_rdydata_s1_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (pio_rdydata_s1_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (pio_rdydata_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_demux_001_src12_ready),                                                      //              cp.ready
		.cp_valid                (cmd_xbar_demux_001_src12_valid),                                                      //                .valid
		.cp_data                 (cmd_xbar_demux_001_src12_data),                                                       //                .data
		.cp_startofpacket        (cmd_xbar_demux_001_src12_startofpacket),                                              //                .startofpacket
		.cp_endofpacket          (cmd_xbar_demux_001_src12_endofpacket),                                                //                .endofpacket
		.cp_channel              (cmd_xbar_demux_001_src12_channel),                                                    //                .channel
		.rf_sink_ready           (pio_rdydata_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (pio_rdydata_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (pio_rdydata_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (pio_rdydata_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (pio_rdydata_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (pio_rdydata_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (pio_rdydata_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (pio_rdydata_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (pio_rdydata_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (pio_rdydata_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (pio_rdydata_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (pio_rdydata_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (pio_rdydata_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (pio_rdydata_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (pio_rdydata_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (pio_rdydata_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data)         //                .data
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (77),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) pio_rdydata_s1_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clk_clk),                                                                             //       clk.clk
		.reset             (rst_controller_reset_out_reset),                                                      // clk_reset.reset
		.in_data           (pio_rdydata_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (pio_rdydata_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (pio_rdydata_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (pio_rdydata_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (pio_rdydata_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (pio_rdydata_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (pio_rdydata_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (pio_rdydata_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (pio_rdydata_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (pio_rdydata_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                               // (terminated)
		.csr_read          (1'b0),                                                                                // (terminated)
		.csr_write         (1'b0),                                                                                // (terminated)
		.csr_readdata      (),                                                                                    // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                // (terminated)
		.almost_full_data  (),                                                                                    // (terminated)
		.almost_empty_data (),                                                                                    // (terminated)
		.in_empty          (1'b0),                                                                                // (terminated)
		.out_empty         (),                                                                                    // (terminated)
		.in_error          (1'b0),                                                                                // (terminated)
		.out_error         (),                                                                                    // (terminated)
		.in_channel        (1'b0),                                                                                // (terminated)
		.out_channel       ()                                                                                     // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (66),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (54),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (55),
		.PKT_TRANS_POSTED          (56),
		.PKT_TRANS_WRITE           (57),
		.PKT_TRANS_READ            (58),
		.PKT_TRANS_LOCK            (59),
		.PKT_SRC_ID_H              (70),
		.PKT_SRC_ID_L              (67),
		.PKT_DEST_ID_H             (74),
		.PKT_DEST_ID_L             (71),
		.PKT_BURSTWRAP_H           (65),
		.PKT_BURSTWRAP_L           (63),
		.PKT_BYTE_CNT_H            (62),
		.PKT_BYTE_CNT_L            (60),
		.PKT_PROTECTION_H          (75),
		.PKT_PROTECTION_L          (75),
		.ST_CHANNEL_W              (14),
		.ST_DATA_W                 (76),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1)
	) jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent (
		.clk                     (clk_clk),                                                                                          //             clk.clk
		.reset                   (rst_controller_reset_out_reset),                                                                   //       clk_reset.reset
		.m0_address              (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_demux_001_src2_ready),                                                                    //              cp.ready
		.cp_valid                (cmd_xbar_demux_001_src2_valid),                                                                    //                .valid
		.cp_data                 (cmd_xbar_demux_001_src2_data),                                                                     //                .data
		.cp_startofpacket        (cmd_xbar_demux_001_src2_startofpacket),                                                            //                .startofpacket
		.cp_endofpacket          (cmd_xbar_demux_001_src2_endofpacket),                                                              //                .endofpacket
		.cp_channel              (cmd_xbar_demux_001_src2_channel),                                                                  //                .channel
		.rf_sink_ready           (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data)         //                .data
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (77),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clk_clk),                                                                                          //       clk.clk
		.reset             (rst_controller_reset_out_reset),                                                                   // clk_reset.reset
		.in_data           (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                            // (terminated)
		.csr_read          (1'b0),                                                                                             // (terminated)
		.csr_write         (1'b0),                                                                                             // (terminated)
		.csr_readdata      (),                                                                                                 // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                             // (terminated)
		.almost_full_data  (),                                                                                                 // (terminated)
		.almost_empty_data (),                                                                                                 // (terminated)
		.in_empty          (1'b0),                                                                                             // (terminated)
		.out_empty         (),                                                                                                 // (terminated)
		.in_error          (1'b0),                                                                                             // (terminated)
		.out_error         (),                                                                                                 // (terminated)
		.in_channel        (1'b0),                                                                                             // (terminated)
		.out_channel       ()                                                                                                  // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (66),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (54),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (55),
		.PKT_TRANS_POSTED          (56),
		.PKT_TRANS_WRITE           (57),
		.PKT_TRANS_READ            (58),
		.PKT_TRANS_LOCK            (59),
		.PKT_SRC_ID_H              (70),
		.PKT_SRC_ID_L              (67),
		.PKT_DEST_ID_H             (74),
		.PKT_DEST_ID_L             (71),
		.PKT_BURSTWRAP_H           (65),
		.PKT_BURSTWRAP_L           (63),
		.PKT_BYTE_CNT_H            (62),
		.PKT_BYTE_CNT_L            (60),
		.PKT_PROTECTION_H          (75),
		.PKT_PROTECTION_L          (75),
		.ST_CHANNEL_W              (14),
		.ST_DATA_W                 (76),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1)
	) lcd_control_slave_translator_avalon_universal_slave_0_agent (
		.clk                     (clk_clk),                                                                                //             clk.clk
		.reset                   (rst_controller_reset_out_reset),                                                         //       clk_reset.reset
		.m0_address              (lcd_control_slave_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (lcd_control_slave_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (lcd_control_slave_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (lcd_control_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (lcd_control_slave_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (lcd_control_slave_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (lcd_control_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (lcd_control_slave_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (lcd_control_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (lcd_control_slave_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (lcd_control_slave_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (lcd_control_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (lcd_control_slave_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (lcd_control_slave_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (lcd_control_slave_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (lcd_control_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_demux_001_src8_ready),                                                          //              cp.ready
		.cp_valid                (cmd_xbar_demux_001_src8_valid),                                                          //                .valid
		.cp_data                 (cmd_xbar_demux_001_src8_data),                                                           //                .data
		.cp_startofpacket        (cmd_xbar_demux_001_src8_startofpacket),                                                  //                .startofpacket
		.cp_endofpacket          (cmd_xbar_demux_001_src8_endofpacket),                                                    //                .endofpacket
		.cp_channel              (cmd_xbar_demux_001_src8_channel),                                                        //                .channel
		.rf_sink_ready           (lcd_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (lcd_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (lcd_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (lcd_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (lcd_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (lcd_control_slave_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (lcd_control_slave_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (lcd_control_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (lcd_control_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (lcd_control_slave_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (lcd_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (lcd_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (lcd_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (lcd_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (lcd_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (lcd_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data)         //                .data
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (77),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) lcd_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clk_clk),                                                                                //       clk.clk
		.reset             (rst_controller_reset_out_reset),                                                         // clk_reset.reset
		.in_data           (lcd_control_slave_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (lcd_control_slave_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (lcd_control_slave_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (lcd_control_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (lcd_control_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (lcd_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (lcd_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (lcd_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (lcd_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (lcd_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                  // (terminated)
		.csr_read          (1'b0),                                                                                   // (terminated)
		.csr_write         (1'b0),                                                                                   // (terminated)
		.csr_readdata      (),                                                                                       // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                   // (terminated)
		.almost_full_data  (),                                                                                       // (terminated)
		.almost_empty_data (),                                                                                       // (terminated)
		.in_empty          (1'b0),                                                                                   // (terminated)
		.out_empty         (),                                                                                       // (terminated)
		.in_error          (1'b0),                                                                                   // (terminated)
		.out_error         (),                                                                                       // (terminated)
		.in_channel        (1'b0),                                                                                   // (terminated)
		.out_channel       ()                                                                                        // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (66),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (54),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (55),
		.PKT_TRANS_POSTED          (56),
		.PKT_TRANS_WRITE           (57),
		.PKT_TRANS_READ            (58),
		.PKT_TRANS_LOCK            (59),
		.PKT_SRC_ID_H              (70),
		.PKT_SRC_ID_L              (67),
		.PKT_DEST_ID_H             (74),
		.PKT_DEST_ID_L             (71),
		.PKT_BURSTWRAP_H           (65),
		.PKT_BURSTWRAP_L           (63),
		.PKT_BYTE_CNT_H            (62),
		.PKT_BYTE_CNT_L            (60),
		.PKT_PROTECTION_H          (75),
		.PKT_PROTECTION_L          (75),
		.ST_CHANNEL_W              (14),
		.ST_DATA_W                 (76),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1)
	) pio_ledr_s1_translator_avalon_universal_slave_0_agent (
		.clk                     (clk_clk),                                                                          //             clk.clk
		.reset                   (rst_controller_reset_out_reset),                                                   //       clk_reset.reset
		.m0_address              (pio_ledr_s1_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (pio_ledr_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (pio_ledr_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (pio_ledr_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (pio_ledr_s1_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (pio_ledr_s1_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (pio_ledr_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (pio_ledr_s1_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (pio_ledr_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (pio_ledr_s1_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (pio_ledr_s1_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (pio_ledr_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (pio_ledr_s1_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (pio_ledr_s1_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (pio_ledr_s1_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (pio_ledr_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_demux_001_src5_ready),                                                    //              cp.ready
		.cp_valid                (cmd_xbar_demux_001_src5_valid),                                                    //                .valid
		.cp_data                 (cmd_xbar_demux_001_src5_data),                                                     //                .data
		.cp_startofpacket        (cmd_xbar_demux_001_src5_startofpacket),                                            //                .startofpacket
		.cp_endofpacket          (cmd_xbar_demux_001_src5_endofpacket),                                              //                .endofpacket
		.cp_channel              (cmd_xbar_demux_001_src5_channel),                                                  //                .channel
		.rf_sink_ready           (pio_ledr_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (pio_ledr_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (pio_ledr_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (pio_ledr_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (pio_ledr_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (pio_ledr_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (pio_ledr_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (pio_ledr_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (pio_ledr_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (pio_ledr_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (pio_ledr_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (pio_ledr_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (pio_ledr_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (pio_ledr_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (pio_ledr_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (pio_ledr_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data)         //                .data
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (77),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) pio_ledr_s1_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clk_clk),                                                                          //       clk.clk
		.reset             (rst_controller_reset_out_reset),                                                   // clk_reset.reset
		.in_data           (pio_ledr_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (pio_ledr_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (pio_ledr_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (pio_ledr_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (pio_ledr_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (pio_ledr_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (pio_ledr_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (pio_ledr_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (pio_ledr_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (pio_ledr_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                            // (terminated)
		.csr_read          (1'b0),                                                                             // (terminated)
		.csr_write         (1'b0),                                                                             // (terminated)
		.csr_readdata      (),                                                                                 // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                             // (terminated)
		.almost_full_data  (),                                                                                 // (terminated)
		.almost_empty_data (),                                                                                 // (terminated)
		.in_empty          (1'b0),                                                                             // (terminated)
		.out_empty         (),                                                                                 // (terminated)
		.in_error          (1'b0),                                                                             // (terminated)
		.out_error         (),                                                                                 // (terminated)
		.in_channel        (1'b0),                                                                             // (terminated)
		.out_channel       ()                                                                                  // (terminated)
	);

	altera_merlin_master_agent #(
		.PKT_PROTECTION_H          (75),
		.PKT_PROTECTION_L          (75),
		.PKT_BEGIN_BURST           (66),
		.PKT_BURSTWRAP_H           (65),
		.PKT_BURSTWRAP_L           (63),
		.PKT_BYTE_CNT_H            (62),
		.PKT_BYTE_CNT_L            (60),
		.PKT_ADDR_H                (54),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (55),
		.PKT_TRANS_POSTED          (56),
		.PKT_TRANS_WRITE           (57),
		.PKT_TRANS_READ            (58),
		.PKT_TRANS_LOCK            (59),
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_SRC_ID_H              (70),
		.PKT_SRC_ID_L              (67),
		.PKT_DEST_ID_H             (74),
		.PKT_DEST_ID_L             (71),
		.ST_DATA_W                 (76),
		.ST_CHANNEL_W              (14),
		.AV_BURSTCOUNT_W           (3),
		.SUPPRESS_0_BYTEEN_RSP     (0),
		.ID                        (0),
		.BURSTWRAP_VALUE           (3)
	) nios2_qsys_instruction_master_translator_avalon_universal_master_0_agent (
		.clk              (clk_clk),                                                                                   //       clk.clk
		.reset            (rst_controller_reset_out_reset),                                                            // clk_reset.reset
		.av_address       (nios2_qsys_instruction_master_translator_avalon_universal_master_0_address),                //        av.address
		.av_write         (nios2_qsys_instruction_master_translator_avalon_universal_master_0_write),                  //          .write
		.av_read          (nios2_qsys_instruction_master_translator_avalon_universal_master_0_read),                   //          .read
		.av_writedata     (nios2_qsys_instruction_master_translator_avalon_universal_master_0_writedata),              //          .writedata
		.av_readdata      (nios2_qsys_instruction_master_translator_avalon_universal_master_0_readdata),               //          .readdata
		.av_waitrequest   (nios2_qsys_instruction_master_translator_avalon_universal_master_0_waitrequest),            //          .waitrequest
		.av_readdatavalid (nios2_qsys_instruction_master_translator_avalon_universal_master_0_readdatavalid),          //          .readdatavalid
		.av_byteenable    (nios2_qsys_instruction_master_translator_avalon_universal_master_0_byteenable),             //          .byteenable
		.av_burstcount    (nios2_qsys_instruction_master_translator_avalon_universal_master_0_burstcount),             //          .burstcount
		.av_debugaccess   (nios2_qsys_instruction_master_translator_avalon_universal_master_0_debugaccess),            //          .debugaccess
		.av_lock          (nios2_qsys_instruction_master_translator_avalon_universal_master_0_lock),                   //          .lock
		.cp_valid         (nios2_qsys_instruction_master_translator_avalon_universal_master_0_agent_cp_valid),         //        cp.valid
		.cp_data          (nios2_qsys_instruction_master_translator_avalon_universal_master_0_agent_cp_data),          //          .data
		.cp_startofpacket (nios2_qsys_instruction_master_translator_avalon_universal_master_0_agent_cp_startofpacket), //          .startofpacket
		.cp_endofpacket   (nios2_qsys_instruction_master_translator_avalon_universal_master_0_agent_cp_endofpacket),   //          .endofpacket
		.cp_ready         (nios2_qsys_instruction_master_translator_avalon_universal_master_0_agent_cp_ready),         //          .ready
		.rp_valid         (limiter_rsp_src_valid),                                                                     //        rp.valid
		.rp_data          (limiter_rsp_src_data),                                                                      //          .data
		.rp_channel       (limiter_rsp_src_channel),                                                                   //          .channel
		.rp_startofpacket (limiter_rsp_src_startofpacket),                                                             //          .startofpacket
		.rp_endofpacket   (limiter_rsp_src_endofpacket),                                                               //          .endofpacket
		.rp_ready         (limiter_rsp_src_ready)                                                                      //          .ready
	);

	altera_merlin_master_agent #(
		.PKT_PROTECTION_H          (75),
		.PKT_PROTECTION_L          (75),
		.PKT_BEGIN_BURST           (66),
		.PKT_BURSTWRAP_H           (65),
		.PKT_BURSTWRAP_L           (63),
		.PKT_BYTE_CNT_H            (62),
		.PKT_BYTE_CNT_L            (60),
		.PKT_ADDR_H                (54),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (55),
		.PKT_TRANS_POSTED          (56),
		.PKT_TRANS_WRITE           (57),
		.PKT_TRANS_READ            (58),
		.PKT_TRANS_LOCK            (59),
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_SRC_ID_H              (70),
		.PKT_SRC_ID_L              (67),
		.PKT_DEST_ID_H             (74),
		.PKT_DEST_ID_L             (71),
		.ST_DATA_W                 (76),
		.ST_CHANNEL_W              (14),
		.AV_BURSTCOUNT_W           (3),
		.SUPPRESS_0_BYTEEN_RSP     (0),
		.ID                        (1),
		.BURSTWRAP_VALUE           (7)
	) nios2_qsys_data_master_translator_avalon_universal_master_0_agent (
		.clk              (clk_clk),                                                                            //       clk.clk
		.reset            (rst_controller_reset_out_reset),                                                     // clk_reset.reset
		.av_address       (nios2_qsys_data_master_translator_avalon_universal_master_0_address),                //        av.address
		.av_write         (nios2_qsys_data_master_translator_avalon_universal_master_0_write),                  //          .write
		.av_read          (nios2_qsys_data_master_translator_avalon_universal_master_0_read),                   //          .read
		.av_writedata     (nios2_qsys_data_master_translator_avalon_universal_master_0_writedata),              //          .writedata
		.av_readdata      (nios2_qsys_data_master_translator_avalon_universal_master_0_readdata),               //          .readdata
		.av_waitrequest   (nios2_qsys_data_master_translator_avalon_universal_master_0_waitrequest),            //          .waitrequest
		.av_readdatavalid (nios2_qsys_data_master_translator_avalon_universal_master_0_readdatavalid),          //          .readdatavalid
		.av_byteenable    (nios2_qsys_data_master_translator_avalon_universal_master_0_byteenable),             //          .byteenable
		.av_burstcount    (nios2_qsys_data_master_translator_avalon_universal_master_0_burstcount),             //          .burstcount
		.av_debugaccess   (nios2_qsys_data_master_translator_avalon_universal_master_0_debugaccess),            //          .debugaccess
		.av_lock          (nios2_qsys_data_master_translator_avalon_universal_master_0_lock),                   //          .lock
		.cp_valid         (nios2_qsys_data_master_translator_avalon_universal_master_0_agent_cp_valid),         //        cp.valid
		.cp_data          (nios2_qsys_data_master_translator_avalon_universal_master_0_agent_cp_data),          //          .data
		.cp_startofpacket (nios2_qsys_data_master_translator_avalon_universal_master_0_agent_cp_startofpacket), //          .startofpacket
		.cp_endofpacket   (nios2_qsys_data_master_translator_avalon_universal_master_0_agent_cp_endofpacket),   //          .endofpacket
		.cp_ready         (nios2_qsys_data_master_translator_avalon_universal_master_0_agent_cp_ready),         //          .ready
		.rp_valid         (limiter_001_rsp_src_valid),                                                          //        rp.valid
		.rp_data          (limiter_001_rsp_src_data),                                                           //          .data
		.rp_channel       (limiter_001_rsp_src_channel),                                                        //          .channel
		.rp_startofpacket (limiter_001_rsp_src_startofpacket),                                                  //          .startofpacket
		.rp_endofpacket   (limiter_001_rsp_src_endofpacket),                                                    //          .endofpacket
		.rp_ready         (limiter_001_rsp_src_ready)                                                           //          .ready
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (66),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (54),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (55),
		.PKT_TRANS_POSTED          (56),
		.PKT_TRANS_WRITE           (57),
		.PKT_TRANS_READ            (58),
		.PKT_TRANS_LOCK            (59),
		.PKT_SRC_ID_H              (70),
		.PKT_SRC_ID_L              (67),
		.PKT_DEST_ID_H             (74),
		.PKT_DEST_ID_L             (71),
		.PKT_BURSTWRAP_H           (65),
		.PKT_BURSTWRAP_L           (63),
		.PKT_BYTE_CNT_H            (62),
		.PKT_BYTE_CNT_L            (60),
		.PKT_PROTECTION_H          (75),
		.PKT_PROTECTION_L          (75),
		.ST_CHANNEL_W              (14),
		.ST_DATA_W                 (76),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1)
	) onchip_memory_s1_translator_avalon_universal_slave_0_agent (
		.clk                     (clk_clk),                                                                               //             clk.clk
		.reset                   (rst_controller_reset_out_reset),                                                        //       clk_reset.reset
		.m0_address              (onchip_memory_s1_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (onchip_memory_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (onchip_memory_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (onchip_memory_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (onchip_memory_s1_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (onchip_memory_s1_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (onchip_memory_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (onchip_memory_s1_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (onchip_memory_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (onchip_memory_s1_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (onchip_memory_s1_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (onchip_memory_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (onchip_memory_s1_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (onchip_memory_s1_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (onchip_memory_s1_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (onchip_memory_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_mux_001_src_ready),                                                            //              cp.ready
		.cp_valid                (cmd_xbar_mux_001_src_valid),                                                            //                .valid
		.cp_data                 (cmd_xbar_mux_001_src_data),                                                             //                .data
		.cp_startofpacket        (cmd_xbar_mux_001_src_startofpacket),                                                    //                .startofpacket
		.cp_endofpacket          (cmd_xbar_mux_001_src_endofpacket),                                                      //                .endofpacket
		.cp_channel              (cmd_xbar_mux_001_src_channel),                                                          //                .channel
		.rf_sink_ready           (onchip_memory_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (onchip_memory_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (onchip_memory_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (onchip_memory_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (onchip_memory_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (onchip_memory_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (onchip_memory_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (onchip_memory_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (onchip_memory_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (onchip_memory_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (onchip_memory_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (onchip_memory_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (onchip_memory_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (onchip_memory_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (onchip_memory_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (onchip_memory_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data)         //                .data
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (77),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) onchip_memory_s1_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clk_clk),                                                                               //       clk.clk
		.reset             (rst_controller_reset_out_reset),                                                        // clk_reset.reset
		.in_data           (onchip_memory_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (onchip_memory_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (onchip_memory_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (onchip_memory_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (onchip_memory_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (onchip_memory_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (onchip_memory_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (onchip_memory_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (onchip_memory_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (onchip_memory_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                 // (terminated)
		.csr_read          (1'b0),                                                                                  // (terminated)
		.csr_write         (1'b0),                                                                                  // (terminated)
		.csr_readdata      (),                                                                                      // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                  // (terminated)
		.almost_full_data  (),                                                                                      // (terminated)
		.almost_empty_data (),                                                                                      // (terminated)
		.in_empty          (1'b0),                                                                                  // (terminated)
		.out_empty         (),                                                                                      // (terminated)
		.in_error          (1'b0),                                                                                  // (terminated)
		.out_error         (),                                                                                      // (terminated)
		.in_channel        (1'b0),                                                                                  // (terminated)
		.out_channel       ()                                                                                       // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (66),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (54),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (55),
		.PKT_TRANS_POSTED          (56),
		.PKT_TRANS_WRITE           (57),
		.PKT_TRANS_READ            (58),
		.PKT_TRANS_LOCK            (59),
		.PKT_SRC_ID_H              (70),
		.PKT_SRC_ID_L              (67),
		.PKT_DEST_ID_H             (74),
		.PKT_DEST_ID_L             (71),
		.PKT_BURSTWRAP_H           (65),
		.PKT_BURSTWRAP_L           (63),
		.PKT_BYTE_CNT_H            (62),
		.PKT_BYTE_CNT_L            (60),
		.PKT_PROTECTION_H          (75),
		.PKT_PROTECTION_L          (75),
		.ST_CHANNEL_W              (14),
		.ST_DATA_W                 (76),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1)
	) pio_sw_s1_translator_avalon_universal_slave_0_agent (
		.clk                     (clk_clk),                                                                        //             clk.clk
		.reset                   (rst_controller_reset_out_reset),                                                 //       clk_reset.reset
		.m0_address              (pio_sw_s1_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (pio_sw_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (pio_sw_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (pio_sw_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (pio_sw_s1_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (pio_sw_s1_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (pio_sw_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (pio_sw_s1_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (pio_sw_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (pio_sw_s1_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (pio_sw_s1_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (pio_sw_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (pio_sw_s1_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (pio_sw_s1_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (pio_sw_s1_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (pio_sw_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_demux_001_src6_ready),                                                  //              cp.ready
		.cp_valid                (cmd_xbar_demux_001_src6_valid),                                                  //                .valid
		.cp_data                 (cmd_xbar_demux_001_src6_data),                                                   //                .data
		.cp_startofpacket        (cmd_xbar_demux_001_src6_startofpacket),                                          //                .startofpacket
		.cp_endofpacket          (cmd_xbar_demux_001_src6_endofpacket),                                            //                .endofpacket
		.cp_channel              (cmd_xbar_demux_001_src6_channel),                                                //                .channel
		.rf_sink_ready           (pio_sw_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (pio_sw_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (pio_sw_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (pio_sw_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (pio_sw_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (pio_sw_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (pio_sw_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (pio_sw_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (pio_sw_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (pio_sw_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (pio_sw_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (pio_sw_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (pio_sw_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (pio_sw_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (pio_sw_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (pio_sw_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data)         //                .data
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (77),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) pio_sw_s1_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clk_clk),                                                                        //       clk.clk
		.reset             (rst_controller_reset_out_reset),                                                 // clk_reset.reset
		.in_data           (pio_sw_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (pio_sw_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (pio_sw_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (pio_sw_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (pio_sw_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (pio_sw_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (pio_sw_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (pio_sw_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (pio_sw_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (pio_sw_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                          // (terminated)
		.csr_read          (1'b0),                                                                           // (terminated)
		.csr_write         (1'b0),                                                                           // (terminated)
		.csr_readdata      (),                                                                               // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                           // (terminated)
		.almost_full_data  (),                                                                               // (terminated)
		.almost_empty_data (),                                                                               // (terminated)
		.in_empty          (1'b0),                                                                           // (terminated)
		.out_empty         (),                                                                               // (terminated)
		.in_error          (1'b0),                                                                           // (terminated)
		.out_error         (),                                                                               // (terminated)
		.in_channel        (1'b0),                                                                           // (terminated)
		.out_channel       ()                                                                                // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (66),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (54),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (55),
		.PKT_TRANS_POSTED          (56),
		.PKT_TRANS_WRITE           (57),
		.PKT_TRANS_READ            (58),
		.PKT_TRANS_LOCK            (59),
		.PKT_SRC_ID_H              (70),
		.PKT_SRC_ID_L              (67),
		.PKT_DEST_ID_H             (74),
		.PKT_DEST_ID_L             (71),
		.PKT_BURSTWRAP_H           (65),
		.PKT_BURSTWRAP_L           (63),
		.PKT_BYTE_CNT_H            (62),
		.PKT_BYTE_CNT_L            (60),
		.PKT_PROTECTION_H          (75),
		.PKT_PROTECTION_L          (75),
		.ST_CHANNEL_W              (14),
		.ST_DATA_W                 (76),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1)
	) sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent (
		.clk                     (clk_clk),                                                                                       //             clk.clk
		.reset                   (rst_controller_reset_out_reset),                                                                //       clk_reset.reset
		.m0_address              (sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_demux_001_src3_ready),                                                                 //              cp.ready
		.cp_valid                (cmd_xbar_demux_001_src3_valid),                                                                 //                .valid
		.cp_data                 (cmd_xbar_demux_001_src3_data),                                                                  //                .data
		.cp_startofpacket        (cmd_xbar_demux_001_src3_startofpacket),                                                         //                .startofpacket
		.cp_endofpacket          (cmd_xbar_demux_001_src3_endofpacket),                                                           //                .endofpacket
		.cp_channel              (cmd_xbar_demux_001_src3_channel),                                                               //                .channel
		.rf_sink_ready           (sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data)         //                .data
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (77),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clk_clk),                                                                                       //       clk.clk
		.reset             (rst_controller_reset_out_reset),                                                                // clk_reset.reset
		.in_data           (sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                         // (terminated)
		.csr_read          (1'b0),                                                                                          // (terminated)
		.csr_write         (1'b0),                                                                                          // (terminated)
		.csr_readdata      (),                                                                                              // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                          // (terminated)
		.almost_full_data  (),                                                                                              // (terminated)
		.almost_empty_data (),                                                                                              // (terminated)
		.in_empty          (1'b0),                                                                                          // (terminated)
		.out_empty         (),                                                                                              // (terminated)
		.in_error          (1'b0),                                                                                          // (terminated)
		.out_error         (),                                                                                              // (terminated)
		.in_channel        (1'b0),                                                                                          // (terminated)
		.out_channel       ()                                                                                               // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (66),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (54),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (55),
		.PKT_TRANS_POSTED          (56),
		.PKT_TRANS_WRITE           (57),
		.PKT_TRANS_READ            (58),
		.PKT_TRANS_LOCK            (59),
		.PKT_SRC_ID_H              (70),
		.PKT_SRC_ID_L              (67),
		.PKT_DEST_ID_H             (74),
		.PKT_DEST_ID_L             (71),
		.PKT_BURSTWRAP_H           (65),
		.PKT_BURSTWRAP_L           (63),
		.PKT_BYTE_CNT_H            (62),
		.PKT_BYTE_CNT_L            (60),
		.PKT_PROTECTION_H          (75),
		.PKT_PROTECTION_L          (75),
		.ST_CHANNEL_W              (14),
		.ST_DATA_W                 (76),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1)
	) nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent (
		.clk                     (clk_clk),                                                                                           //             clk.clk
		.reset                   (rst_controller_reset_out_reset),                                                                    //       clk_reset.reset
		.m0_address              (nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_mux_src_ready),                                                                            //              cp.ready
		.cp_valid                (cmd_xbar_mux_src_valid),                                                                            //                .valid
		.cp_data                 (cmd_xbar_mux_src_data),                                                                             //                .data
		.cp_startofpacket        (cmd_xbar_mux_src_startofpacket),                                                                    //                .startofpacket
		.cp_endofpacket          (cmd_xbar_mux_src_endofpacket),                                                                      //                .endofpacket
		.cp_channel              (cmd_xbar_mux_src_channel),                                                                          //                .channel
		.rf_sink_ready           (nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data)         //                .data
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (77),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clk_clk),                                                                                           //       clk.clk
		.reset             (rst_controller_reset_out_reset),                                                                    // clk_reset.reset
		.in_data           (nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                             // (terminated)
		.csr_read          (1'b0),                                                                                              // (terminated)
		.csr_write         (1'b0),                                                                                              // (terminated)
		.csr_readdata      (),                                                                                                  // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                              // (terminated)
		.almost_full_data  (),                                                                                                  // (terminated)
		.almost_empty_data (),                                                                                                  // (terminated)
		.in_empty          (1'b0),                                                                                              // (terminated)
		.out_empty         (),                                                                                                  // (terminated)
		.in_error          (1'b0),                                                                                              // (terminated)
		.out_error         (),                                                                                                  // (terminated)
		.in_channel        (1'b0),                                                                                              // (terminated)
		.out_channel       ()                                                                                                   // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (66),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (54),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (55),
		.PKT_TRANS_POSTED          (56),
		.PKT_TRANS_WRITE           (57),
		.PKT_TRANS_READ            (58),
		.PKT_TRANS_LOCK            (59),
		.PKT_SRC_ID_H              (70),
		.PKT_SRC_ID_L              (67),
		.PKT_DEST_ID_H             (74),
		.PKT_DEST_ID_L             (71),
		.PKT_BURSTWRAP_H           (65),
		.PKT_BURSTWRAP_L           (63),
		.PKT_BYTE_CNT_H            (62),
		.PKT_BYTE_CNT_L            (60),
		.PKT_PROTECTION_H          (75),
		.PKT_PROTECTION_L          (75),
		.ST_CHANNEL_W              (14),
		.ST_DATA_W                 (76),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1)
	) pio_ledg_s1_translator_avalon_universal_slave_0_agent (
		.clk                     (clk_clk),                                                                          //             clk.clk
		.reset                   (rst_controller_reset_out_reset),                                                   //       clk_reset.reset
		.m0_address              (pio_ledg_s1_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (pio_ledg_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (pio_ledg_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (pio_ledg_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (pio_ledg_s1_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (pio_ledg_s1_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (pio_ledg_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (pio_ledg_s1_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (pio_ledg_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (pio_ledg_s1_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (pio_ledg_s1_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (pio_ledg_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (pio_ledg_s1_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (pio_ledg_s1_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (pio_ledg_s1_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (pio_ledg_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_demux_001_src4_ready),                                                    //              cp.ready
		.cp_valid                (cmd_xbar_demux_001_src4_valid),                                                    //                .valid
		.cp_data                 (cmd_xbar_demux_001_src4_data),                                                     //                .data
		.cp_startofpacket        (cmd_xbar_demux_001_src4_startofpacket),                                            //                .startofpacket
		.cp_endofpacket          (cmd_xbar_demux_001_src4_endofpacket),                                              //                .endofpacket
		.cp_channel              (cmd_xbar_demux_001_src4_channel),                                                  //                .channel
		.rf_sink_ready           (pio_ledg_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (pio_ledg_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (pio_ledg_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (pio_ledg_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (pio_ledg_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (pio_ledg_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (pio_ledg_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (pio_ledg_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (pio_ledg_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (pio_ledg_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (pio_ledg_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (pio_ledg_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (pio_ledg_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (pio_ledg_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (pio_ledg_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (pio_ledg_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data)         //                .data
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (77),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) pio_ledg_s1_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clk_clk),                                                                          //       clk.clk
		.reset             (rst_controller_reset_out_reset),                                                   // clk_reset.reset
		.in_data           (pio_ledg_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (pio_ledg_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (pio_ledg_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (pio_ledg_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (pio_ledg_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (pio_ledg_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (pio_ledg_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (pio_ledg_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (pio_ledg_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (pio_ledg_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                            // (terminated)
		.csr_read          (1'b0),                                                                             // (terminated)
		.csr_write         (1'b0),                                                                             // (terminated)
		.csr_readdata      (),                                                                                 // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                             // (terminated)
		.almost_full_data  (),                                                                                 // (terminated)
		.almost_empty_data (),                                                                                 // (terminated)
		.in_empty          (1'b0),                                                                             // (terminated)
		.out_empty         (),                                                                                 // (terminated)
		.in_error          (1'b0),                                                                             // (terminated)
		.out_error         (),                                                                                 // (terminated)
		.in_channel        (1'b0),                                                                             // (terminated)
		.out_channel       ()                                                                                  // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (66),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (54),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (55),
		.PKT_TRANS_POSTED          (56),
		.PKT_TRANS_WRITE           (57),
		.PKT_TRANS_READ            (58),
		.PKT_TRANS_LOCK            (59),
		.PKT_SRC_ID_H              (70),
		.PKT_SRC_ID_L              (67),
		.PKT_DEST_ID_H             (74),
		.PKT_DEST_ID_L             (71),
		.PKT_BURSTWRAP_H           (65),
		.PKT_BURSTWRAP_L           (63),
		.PKT_BYTE_CNT_H            (62),
		.PKT_BYTE_CNT_L            (60),
		.PKT_PROTECTION_H          (75),
		.PKT_PROTECTION_L          (75),
		.ST_CHANNEL_W              (14),
		.ST_DATA_W                 (76),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1)
	) pio_data_s1_translator_avalon_universal_slave_0_agent (
		.clk                     (clk_clk),                                                                          //             clk.clk
		.reset                   (rst_controller_reset_out_reset),                                                   //       clk_reset.reset
		.m0_address              (pio_data_s1_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (pio_data_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (pio_data_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (pio_data_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (pio_data_s1_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (pio_data_s1_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (pio_data_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (pio_data_s1_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (pio_data_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (pio_data_s1_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (pio_data_s1_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (pio_data_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (pio_data_s1_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (pio_data_s1_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (pio_data_s1_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (pio_data_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_demux_001_src11_ready),                                                   //              cp.ready
		.cp_valid                (cmd_xbar_demux_001_src11_valid),                                                   //                .valid
		.cp_data                 (cmd_xbar_demux_001_src11_data),                                                    //                .data
		.cp_startofpacket        (cmd_xbar_demux_001_src11_startofpacket),                                           //                .startofpacket
		.cp_endofpacket          (cmd_xbar_demux_001_src11_endofpacket),                                             //                .endofpacket
		.cp_channel              (cmd_xbar_demux_001_src11_channel),                                                 //                .channel
		.rf_sink_ready           (pio_data_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (pio_data_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (pio_data_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (pio_data_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (pio_data_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (pio_data_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (pio_data_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (pio_data_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (pio_data_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (pio_data_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (pio_data_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (pio_data_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (pio_data_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (pio_data_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (pio_data_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (pio_data_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data)         //                .data
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (77),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) pio_data_s1_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clk_clk),                                                                          //       clk.clk
		.reset             (rst_controller_reset_out_reset),                                                   // clk_reset.reset
		.in_data           (pio_data_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (pio_data_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (pio_data_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (pio_data_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (pio_data_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (pio_data_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (pio_data_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (pio_data_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (pio_data_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (pio_data_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                            // (terminated)
		.csr_read          (1'b0),                                                                             // (terminated)
		.csr_write         (1'b0),                                                                             // (terminated)
		.csr_readdata      (),                                                                                 // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                             // (terminated)
		.almost_full_data  (),                                                                                 // (terminated)
		.almost_empty_data (),                                                                                 // (terminated)
		.in_empty          (1'b0),                                                                             // (terminated)
		.out_empty         (),                                                                                 // (terminated)
		.in_error          (1'b0),                                                                             // (terminated)
		.out_error         (),                                                                                 // (terminated)
		.in_channel        (1'b0),                                                                             // (terminated)
		.out_channel       ()                                                                                  // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (66),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (54),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (55),
		.PKT_TRANS_POSTED          (56),
		.PKT_TRANS_WRITE           (57),
		.PKT_TRANS_READ            (58),
		.PKT_TRANS_LOCK            (59),
		.PKT_SRC_ID_H              (70),
		.PKT_SRC_ID_L              (67),
		.PKT_DEST_ID_H             (74),
		.PKT_DEST_ID_L             (71),
		.PKT_BURSTWRAP_H           (65),
		.PKT_BURSTWRAP_L           (63),
		.PKT_BYTE_CNT_H            (62),
		.PKT_BYTE_CNT_L            (60),
		.PKT_PROTECTION_H          (75),
		.PKT_PROTECTION_L          (75),
		.ST_CHANNEL_W              (14),
		.ST_DATA_W                 (76),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1)
	) pio_button_s1_translator_avalon_universal_slave_0_agent (
		.clk                     (clk_clk),                                                                            //             clk.clk
		.reset                   (rst_controller_reset_out_reset),                                                     //       clk_reset.reset
		.m0_address              (pio_button_s1_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (pio_button_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (pio_button_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (pio_button_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (pio_button_s1_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (pio_button_s1_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (pio_button_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (pio_button_s1_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (pio_button_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (pio_button_s1_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (pio_button_s1_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (pio_button_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (pio_button_s1_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (pio_button_s1_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (pio_button_s1_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (pio_button_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_demux_001_src7_ready),                                                      //              cp.ready
		.cp_valid                (cmd_xbar_demux_001_src7_valid),                                                      //                .valid
		.cp_data                 (cmd_xbar_demux_001_src7_data),                                                       //                .data
		.cp_startofpacket        (cmd_xbar_demux_001_src7_startofpacket),                                              //                .startofpacket
		.cp_endofpacket          (cmd_xbar_demux_001_src7_endofpacket),                                                //                .endofpacket
		.cp_channel              (cmd_xbar_demux_001_src7_channel),                                                    //                .channel
		.rf_sink_ready           (pio_button_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (pio_button_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (pio_button_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (pio_button_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (pio_button_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (pio_button_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (pio_button_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (pio_button_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (pio_button_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (pio_button_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (pio_button_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (pio_button_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (pio_button_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (pio_button_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (pio_button_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (pio_button_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data)         //                .data
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (77),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) pio_button_s1_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clk_clk),                                                                            //       clk.clk
		.reset             (rst_controller_reset_out_reset),                                                     // clk_reset.reset
		.in_data           (pio_button_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (pio_button_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (pio_button_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (pio_button_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (pio_button_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (pio_button_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (pio_button_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (pio_button_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (pio_button_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (pio_button_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                              // (terminated)
		.csr_read          (1'b0),                                                                               // (terminated)
		.csr_write         (1'b0),                                                                               // (terminated)
		.csr_readdata      (),                                                                                   // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                               // (terminated)
		.almost_full_data  (),                                                                                   // (terminated)
		.almost_empty_data (),                                                                                   // (terminated)
		.in_empty          (1'b0),                                                                               // (terminated)
		.out_empty         (),                                                                                   // (terminated)
		.in_error          (1'b0),                                                                               // (terminated)
		.out_error         (),                                                                                   // (terminated)
		.in_channel        (1'b0),                                                                               // (terminated)
		.out_channel       ()                                                                                    // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (66),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (54),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (55),
		.PKT_TRANS_POSTED          (56),
		.PKT_TRANS_WRITE           (57),
		.PKT_TRANS_READ            (58),
		.PKT_TRANS_LOCK            (59),
		.PKT_SRC_ID_H              (70),
		.PKT_SRC_ID_L              (67),
		.PKT_DEST_ID_H             (74),
		.PKT_DEST_ID_L             (71),
		.PKT_BURSTWRAP_H           (65),
		.PKT_BURSTWRAP_L           (63),
		.PKT_BYTE_CNT_H            (62),
		.PKT_BYTE_CNT_L            (60),
		.PKT_PROTECTION_H          (75),
		.PKT_PROTECTION_L          (75),
		.ST_CHANNEL_W              (14),
		.ST_DATA_W                 (76),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1)
	) timer_0_s1_translator_avalon_universal_slave_0_agent (
		.clk                     (clk_clk),                                                                         //             clk.clk
		.reset                   (rst_controller_reset_out_reset),                                                  //       clk_reset.reset
		.m0_address              (timer_0_s1_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (timer_0_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (timer_0_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (timer_0_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (timer_0_s1_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (timer_0_s1_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (timer_0_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (timer_0_s1_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (timer_0_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (timer_0_s1_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (timer_0_s1_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (timer_0_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (timer_0_s1_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (timer_0_s1_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (timer_0_s1_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (timer_0_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_demux_001_src10_ready),                                                  //              cp.ready
		.cp_valid                (cmd_xbar_demux_001_src10_valid),                                                  //                .valid
		.cp_data                 (cmd_xbar_demux_001_src10_data),                                                   //                .data
		.cp_startofpacket        (cmd_xbar_demux_001_src10_startofpacket),                                          //                .startofpacket
		.cp_endofpacket          (cmd_xbar_demux_001_src10_endofpacket),                                            //                .endofpacket
		.cp_channel              (cmd_xbar_demux_001_src10_channel),                                                //                .channel
		.rf_sink_ready           (timer_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (timer_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (timer_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (timer_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (timer_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (timer_0_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (timer_0_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (timer_0_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (timer_0_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (timer_0_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (timer_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (timer_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (timer_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (timer_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (timer_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (timer_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data)         //                .data
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (77),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) timer_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clk_clk),                                                                         //       clk.clk
		.reset             (rst_controller_reset_out_reset),                                                  // clk_reset.reset
		.in_data           (timer_0_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (timer_0_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (timer_0_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (timer_0_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (timer_0_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (timer_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (timer_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (timer_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (timer_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (timer_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                           // (terminated)
		.csr_read          (1'b0),                                                                            // (terminated)
		.csr_write         (1'b0),                                                                            // (terminated)
		.csr_readdata      (),                                                                                // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                            // (terminated)
		.almost_full_data  (),                                                                                // (terminated)
		.almost_empty_data (),                                                                                // (terminated)
		.in_empty          (1'b0),                                                                            // (terminated)
		.out_empty         (),                                                                                // (terminated)
		.in_error          (1'b0),                                                                            // (terminated)
		.out_error         (),                                                                                // (terminated)
		.in_channel        (1'b0),                                                                            // (terminated)
		.out_channel       ()                                                                                 // (terminated)
	);

	Nios1_addr_router addr_router (
		.sink_ready         (nios2_qsys_instruction_master_translator_avalon_universal_master_0_agent_cp_ready),         //      sink.ready
		.sink_valid         (nios2_qsys_instruction_master_translator_avalon_universal_master_0_agent_cp_valid),         //          .valid
		.sink_data          (nios2_qsys_instruction_master_translator_avalon_universal_master_0_agent_cp_data),          //          .data
		.sink_startofpacket (nios2_qsys_instruction_master_translator_avalon_universal_master_0_agent_cp_startofpacket), //          .startofpacket
		.sink_endofpacket   (nios2_qsys_instruction_master_translator_avalon_universal_master_0_agent_cp_endofpacket),   //          .endofpacket
		.clk                (clk_clk),                                                                                   //       clk.clk
		.reset              (rst_controller_reset_out_reset),                                                            // clk_reset.reset
		.src_ready          (addr_router_src_ready),                                                                     //       src.ready
		.src_valid          (addr_router_src_valid),                                                                     //          .valid
		.src_data           (addr_router_src_data),                                                                      //          .data
		.src_channel        (addr_router_src_channel),                                                                   //          .channel
		.src_startofpacket  (addr_router_src_startofpacket),                                                             //          .startofpacket
		.src_endofpacket    (addr_router_src_endofpacket)                                                                //          .endofpacket
	);

	Nios1_addr_router_001 addr_router_001 (
		.sink_ready         (nios2_qsys_data_master_translator_avalon_universal_master_0_agent_cp_ready),         //      sink.ready
		.sink_valid         (nios2_qsys_data_master_translator_avalon_universal_master_0_agent_cp_valid),         //          .valid
		.sink_data          (nios2_qsys_data_master_translator_avalon_universal_master_0_agent_cp_data),          //          .data
		.sink_startofpacket (nios2_qsys_data_master_translator_avalon_universal_master_0_agent_cp_startofpacket), //          .startofpacket
		.sink_endofpacket   (nios2_qsys_data_master_translator_avalon_universal_master_0_agent_cp_endofpacket),   //          .endofpacket
		.clk                (clk_clk),                                                                            //       clk.clk
		.reset              (rst_controller_reset_out_reset),                                                     // clk_reset.reset
		.src_ready          (addr_router_001_src_ready),                                                          //       src.ready
		.src_valid          (addr_router_001_src_valid),                                                          //          .valid
		.src_data           (addr_router_001_src_data),                                                           //          .data
		.src_channel        (addr_router_001_src_channel),                                                        //          .channel
		.src_startofpacket  (addr_router_001_src_startofpacket),                                                  //          .startofpacket
		.src_endofpacket    (addr_router_001_src_endofpacket)                                                     //          .endofpacket
	);

	Nios1_id_router id_router (
		.sink_ready         (nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (clk_clk),                                                                                 //       clk.clk
		.reset              (rst_controller_reset_out_reset),                                                          // clk_reset.reset
		.src_ready          (id_router_src_ready),                                                                     //       src.ready
		.src_valid          (id_router_src_valid),                                                                     //          .valid
		.src_data           (id_router_src_data),                                                                      //          .data
		.src_channel        (id_router_src_channel),                                                                   //          .channel
		.src_startofpacket  (id_router_src_startofpacket),                                                             //          .startofpacket
		.src_endofpacket    (id_router_src_endofpacket)                                                                //          .endofpacket
	);

	Nios1_id_router id_router_001 (
		.sink_ready         (onchip_memory_s1_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (onchip_memory_s1_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (onchip_memory_s1_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (onchip_memory_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (onchip_memory_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (clk_clk),                                                                     //       clk.clk
		.reset              (rst_controller_reset_out_reset),                                              // clk_reset.reset
		.src_ready          (id_router_001_src_ready),                                                     //       src.ready
		.src_valid          (id_router_001_src_valid),                                                     //          .valid
		.src_data           (id_router_001_src_data),                                                      //          .data
		.src_channel        (id_router_001_src_channel),                                                   //          .channel
		.src_startofpacket  (id_router_001_src_startofpacket),                                             //          .startofpacket
		.src_endofpacket    (id_router_001_src_endofpacket)                                                //          .endofpacket
	);

	Nios1_id_router_002 id_router_002 (
		.sink_ready         (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (clk_clk),                                                                                //       clk.clk
		.reset              (rst_controller_reset_out_reset),                                                         // clk_reset.reset
		.src_ready          (id_router_002_src_ready),                                                                //       src.ready
		.src_valid          (id_router_002_src_valid),                                                                //          .valid
		.src_data           (id_router_002_src_data),                                                                 //          .data
		.src_channel        (id_router_002_src_channel),                                                              //          .channel
		.src_startofpacket  (id_router_002_src_startofpacket),                                                        //          .startofpacket
		.src_endofpacket    (id_router_002_src_endofpacket)                                                           //          .endofpacket
	);

	Nios1_id_router_002 id_router_003 (
		.sink_ready         (sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (clk_clk),                                                                             //       clk.clk
		.reset              (rst_controller_reset_out_reset),                                                      // clk_reset.reset
		.src_ready          (id_router_003_src_ready),                                                             //       src.ready
		.src_valid          (id_router_003_src_valid),                                                             //          .valid
		.src_data           (id_router_003_src_data),                                                              //          .data
		.src_channel        (id_router_003_src_channel),                                                           //          .channel
		.src_startofpacket  (id_router_003_src_startofpacket),                                                     //          .startofpacket
		.src_endofpacket    (id_router_003_src_endofpacket)                                                        //          .endofpacket
	);

	Nios1_id_router_002 id_router_004 (
		.sink_ready         (pio_ledg_s1_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (pio_ledg_s1_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (pio_ledg_s1_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (pio_ledg_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (pio_ledg_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (clk_clk),                                                                //       clk.clk
		.reset              (rst_controller_reset_out_reset),                                         // clk_reset.reset
		.src_ready          (id_router_004_src_ready),                                                //       src.ready
		.src_valid          (id_router_004_src_valid),                                                //          .valid
		.src_data           (id_router_004_src_data),                                                 //          .data
		.src_channel        (id_router_004_src_channel),                                              //          .channel
		.src_startofpacket  (id_router_004_src_startofpacket),                                        //          .startofpacket
		.src_endofpacket    (id_router_004_src_endofpacket)                                           //          .endofpacket
	);

	Nios1_id_router_002 id_router_005 (
		.sink_ready         (pio_ledr_s1_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (pio_ledr_s1_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (pio_ledr_s1_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (pio_ledr_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (pio_ledr_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (clk_clk),                                                                //       clk.clk
		.reset              (rst_controller_reset_out_reset),                                         // clk_reset.reset
		.src_ready          (id_router_005_src_ready),                                                //       src.ready
		.src_valid          (id_router_005_src_valid),                                                //          .valid
		.src_data           (id_router_005_src_data),                                                 //          .data
		.src_channel        (id_router_005_src_channel),                                              //          .channel
		.src_startofpacket  (id_router_005_src_startofpacket),                                        //          .startofpacket
		.src_endofpacket    (id_router_005_src_endofpacket)                                           //          .endofpacket
	);

	Nios1_id_router_002 id_router_006 (
		.sink_ready         (pio_sw_s1_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (pio_sw_s1_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (pio_sw_s1_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (pio_sw_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (pio_sw_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (clk_clk),                                                              //       clk.clk
		.reset              (rst_controller_reset_out_reset),                                       // clk_reset.reset
		.src_ready          (id_router_006_src_ready),                                              //       src.ready
		.src_valid          (id_router_006_src_valid),                                              //          .valid
		.src_data           (id_router_006_src_data),                                               //          .data
		.src_channel        (id_router_006_src_channel),                                            //          .channel
		.src_startofpacket  (id_router_006_src_startofpacket),                                      //          .startofpacket
		.src_endofpacket    (id_router_006_src_endofpacket)                                         //          .endofpacket
	);

	Nios1_id_router_002 id_router_007 (
		.sink_ready         (pio_button_s1_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (pio_button_s1_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (pio_button_s1_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (pio_button_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (pio_button_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (clk_clk),                                                                  //       clk.clk
		.reset              (rst_controller_reset_out_reset),                                           // clk_reset.reset
		.src_ready          (id_router_007_src_ready),                                                  //       src.ready
		.src_valid          (id_router_007_src_valid),                                                  //          .valid
		.src_data           (id_router_007_src_data),                                                   //          .data
		.src_channel        (id_router_007_src_channel),                                                //          .channel
		.src_startofpacket  (id_router_007_src_startofpacket),                                          //          .startofpacket
		.src_endofpacket    (id_router_007_src_endofpacket)                                             //          .endofpacket
	);

	Nios1_id_router_002 id_router_008 (
		.sink_ready         (lcd_control_slave_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (lcd_control_slave_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (lcd_control_slave_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (lcd_control_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (lcd_control_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (clk_clk),                                                                      //       clk.clk
		.reset              (rst_controller_reset_out_reset),                                               // clk_reset.reset
		.src_ready          (id_router_008_src_ready),                                                      //       src.ready
		.src_valid          (id_router_008_src_valid),                                                      //          .valid
		.src_data           (id_router_008_src_data),                                                       //          .data
		.src_channel        (id_router_008_src_channel),                                                    //          .channel
		.src_startofpacket  (id_router_008_src_startofpacket),                                              //          .startofpacket
		.src_endofpacket    (id_router_008_src_endofpacket)                                                 //          .endofpacket
	);

	Nios1_id_router_002 id_router_009 (
		.sink_ready         (uart_s1_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (uart_s1_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (uart_s1_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (uart_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (uart_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (clk_clk),                                                            //       clk.clk
		.reset              (rst_controller_reset_out_reset),                                     // clk_reset.reset
		.src_ready          (id_router_009_src_ready),                                            //       src.ready
		.src_valid          (id_router_009_src_valid),                                            //          .valid
		.src_data           (id_router_009_src_data),                                             //          .data
		.src_channel        (id_router_009_src_channel),                                          //          .channel
		.src_startofpacket  (id_router_009_src_startofpacket),                                    //          .startofpacket
		.src_endofpacket    (id_router_009_src_endofpacket)                                       //          .endofpacket
	);

	Nios1_id_router_002 id_router_010 (
		.sink_ready         (timer_0_s1_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (timer_0_s1_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (timer_0_s1_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (timer_0_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (timer_0_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (clk_clk),                                                               //       clk.clk
		.reset              (rst_controller_reset_out_reset),                                        // clk_reset.reset
		.src_ready          (id_router_010_src_ready),                                               //       src.ready
		.src_valid          (id_router_010_src_valid),                                               //          .valid
		.src_data           (id_router_010_src_data),                                                //          .data
		.src_channel        (id_router_010_src_channel),                                             //          .channel
		.src_startofpacket  (id_router_010_src_startofpacket),                                       //          .startofpacket
		.src_endofpacket    (id_router_010_src_endofpacket)                                          //          .endofpacket
	);

	Nios1_id_router_002 id_router_011 (
		.sink_ready         (pio_data_s1_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (pio_data_s1_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (pio_data_s1_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (pio_data_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (pio_data_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (clk_clk),                                                                //       clk.clk
		.reset              (rst_controller_reset_out_reset),                                         // clk_reset.reset
		.src_ready          (id_router_011_src_ready),                                                //       src.ready
		.src_valid          (id_router_011_src_valid),                                                //          .valid
		.src_data           (id_router_011_src_data),                                                 //          .data
		.src_channel        (id_router_011_src_channel),                                              //          .channel
		.src_startofpacket  (id_router_011_src_startofpacket),                                        //          .startofpacket
		.src_endofpacket    (id_router_011_src_endofpacket)                                           //          .endofpacket
	);

	Nios1_id_router_002 id_router_012 (
		.sink_ready         (pio_rdydata_s1_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (pio_rdydata_s1_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (pio_rdydata_s1_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (pio_rdydata_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (pio_rdydata_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (clk_clk),                                                                   //       clk.clk
		.reset              (rst_controller_reset_out_reset),                                            // clk_reset.reset
		.src_ready          (id_router_012_src_ready),                                                   //       src.ready
		.src_valid          (id_router_012_src_valid),                                                   //          .valid
		.src_data           (id_router_012_src_data),                                                    //          .data
		.src_channel        (id_router_012_src_channel),                                                 //          .channel
		.src_startofpacket  (id_router_012_src_startofpacket),                                           //          .startofpacket
		.src_endofpacket    (id_router_012_src_endofpacket)                                              //          .endofpacket
	);

	Nios1_id_router_002 id_router_013 (
		.sink_ready         (pio_dataread_s1_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (pio_dataread_s1_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (pio_dataread_s1_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (pio_dataread_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (pio_dataread_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (clk_clk),                                                                    //       clk.clk
		.reset              (rst_controller_reset_out_reset),                                             // clk_reset.reset
		.src_ready          (id_router_013_src_ready),                                                    //       src.ready
		.src_valid          (id_router_013_src_valid),                                                    //          .valid
		.src_data           (id_router_013_src_data),                                                     //          .data
		.src_channel        (id_router_013_src_channel),                                                  //          .channel
		.src_startofpacket  (id_router_013_src_startofpacket),                                            //          .startofpacket
		.src_endofpacket    (id_router_013_src_endofpacket)                                               //          .endofpacket
	);

	altera_merlin_traffic_limiter #(
		.PKT_DEST_ID_H             (74),
		.PKT_DEST_ID_L             (71),
		.PKT_TRANS_POSTED          (56),
		.MAX_OUTSTANDING_RESPONSES (1),
		.PIPELINED                 (0),
		.ST_DATA_W                 (76),
		.ST_CHANNEL_W              (14),
		.VALID_WIDTH               (14),
		.ENFORCE_ORDER             (1),
		.PKT_BYTE_CNT_H            (62),
		.PKT_BYTE_CNT_L            (60),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32)
	) limiter (
		.clk                    (clk_clk),                        //       clk.clk
		.reset                  (rst_controller_reset_out_reset), // clk_reset.reset
		.cmd_sink_ready         (addr_router_src_ready),          //  cmd_sink.ready
		.cmd_sink_valid         (addr_router_src_valid),          //          .valid
		.cmd_sink_data          (addr_router_src_data),           //          .data
		.cmd_sink_channel       (addr_router_src_channel),        //          .channel
		.cmd_sink_startofpacket (addr_router_src_startofpacket),  //          .startofpacket
		.cmd_sink_endofpacket   (addr_router_src_endofpacket),    //          .endofpacket
		.cmd_src_ready          (limiter_cmd_src_ready),          //   cmd_src.ready
		.cmd_src_data           (limiter_cmd_src_data),           //          .data
		.cmd_src_channel        (limiter_cmd_src_channel),        //          .channel
		.cmd_src_startofpacket  (limiter_cmd_src_startofpacket),  //          .startofpacket
		.cmd_src_endofpacket    (limiter_cmd_src_endofpacket),    //          .endofpacket
		.rsp_sink_ready         (rsp_xbar_mux_src_ready),         //  rsp_sink.ready
		.rsp_sink_valid         (rsp_xbar_mux_src_valid),         //          .valid
		.rsp_sink_channel       (rsp_xbar_mux_src_channel),       //          .channel
		.rsp_sink_data          (rsp_xbar_mux_src_data),          //          .data
		.rsp_sink_startofpacket (rsp_xbar_mux_src_startofpacket), //          .startofpacket
		.rsp_sink_endofpacket   (rsp_xbar_mux_src_endofpacket),   //          .endofpacket
		.rsp_src_ready          (limiter_rsp_src_ready),          //   rsp_src.ready
		.rsp_src_valid          (limiter_rsp_src_valid),          //          .valid
		.rsp_src_data           (limiter_rsp_src_data),           //          .data
		.rsp_src_channel        (limiter_rsp_src_channel),        //          .channel
		.rsp_src_startofpacket  (limiter_rsp_src_startofpacket),  //          .startofpacket
		.rsp_src_endofpacket    (limiter_rsp_src_endofpacket),    //          .endofpacket
		.cmd_src_valid          (limiter_cmd_valid_data)          // cmd_valid.data
	);

	altera_merlin_traffic_limiter #(
		.PKT_DEST_ID_H             (74),
		.PKT_DEST_ID_L             (71),
		.PKT_TRANS_POSTED          (56),
		.MAX_OUTSTANDING_RESPONSES (1),
		.PIPELINED                 (0),
		.ST_DATA_W                 (76),
		.ST_CHANNEL_W              (14),
		.VALID_WIDTH               (14),
		.ENFORCE_ORDER             (1),
		.PKT_BYTE_CNT_H            (62),
		.PKT_BYTE_CNT_L            (60),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32)
	) limiter_001 (
		.clk                    (clk_clk),                            //       clk.clk
		.reset                  (rst_controller_reset_out_reset),     // clk_reset.reset
		.cmd_sink_ready         (addr_router_001_src_ready),          //  cmd_sink.ready
		.cmd_sink_valid         (addr_router_001_src_valid),          //          .valid
		.cmd_sink_data          (addr_router_001_src_data),           //          .data
		.cmd_sink_channel       (addr_router_001_src_channel),        //          .channel
		.cmd_sink_startofpacket (addr_router_001_src_startofpacket),  //          .startofpacket
		.cmd_sink_endofpacket   (addr_router_001_src_endofpacket),    //          .endofpacket
		.cmd_src_ready          (limiter_001_cmd_src_ready),          //   cmd_src.ready
		.cmd_src_data           (limiter_001_cmd_src_data),           //          .data
		.cmd_src_channel        (limiter_001_cmd_src_channel),        //          .channel
		.cmd_src_startofpacket  (limiter_001_cmd_src_startofpacket),  //          .startofpacket
		.cmd_src_endofpacket    (limiter_001_cmd_src_endofpacket),    //          .endofpacket
		.rsp_sink_ready         (rsp_xbar_mux_001_src_ready),         //  rsp_sink.ready
		.rsp_sink_valid         (rsp_xbar_mux_001_src_valid),         //          .valid
		.rsp_sink_channel       (rsp_xbar_mux_001_src_channel),       //          .channel
		.rsp_sink_data          (rsp_xbar_mux_001_src_data),          //          .data
		.rsp_sink_startofpacket (rsp_xbar_mux_001_src_startofpacket), //          .startofpacket
		.rsp_sink_endofpacket   (rsp_xbar_mux_001_src_endofpacket),   //          .endofpacket
		.rsp_src_ready          (limiter_001_rsp_src_ready),          //   rsp_src.ready
		.rsp_src_valid          (limiter_001_rsp_src_valid),          //          .valid
		.rsp_src_data           (limiter_001_rsp_src_data),           //          .data
		.rsp_src_channel        (limiter_001_rsp_src_channel),        //          .channel
		.rsp_src_startofpacket  (limiter_001_rsp_src_startofpacket),  //          .startofpacket
		.rsp_src_endofpacket    (limiter_001_rsp_src_endofpacket),    //          .endofpacket
		.cmd_src_valid          (limiter_001_cmd_valid_data)          // cmd_valid.data
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS        (1),
		.OUTPUT_RESET_SYNC_EDGES ("deassert"),
		.SYNC_DEPTH              (2)
	) rst_controller (
		.reset_in0  (~reset_reset_n),                 // reset_in0.reset
		.clk        (clk_clk),                        //       clk.clk
		.reset_out  (rst_controller_reset_out_reset), // reset_out.reset
		.reset_in1  (1'b0),                           // (terminated)
		.reset_in2  (1'b0),                           // (terminated)
		.reset_in3  (1'b0),                           // (terminated)
		.reset_in4  (1'b0),                           // (terminated)
		.reset_in5  (1'b0),                           // (terminated)
		.reset_in6  (1'b0),                           // (terminated)
		.reset_in7  (1'b0),                           // (terminated)
		.reset_in8  (1'b0),                           // (terminated)
		.reset_in9  (1'b0),                           // (terminated)
		.reset_in10 (1'b0),                           // (terminated)
		.reset_in11 (1'b0),                           // (terminated)
		.reset_in12 (1'b0),                           // (terminated)
		.reset_in13 (1'b0),                           // (terminated)
		.reset_in14 (1'b0),                           // (terminated)
		.reset_in15 (1'b0)                            // (terminated)
	);

	Nios1_cmd_xbar_demux cmd_xbar_demux (
		.clk                (clk_clk),                           //        clk.clk
		.reset              (rst_controller_reset_out_reset),    //  clk_reset.reset
		.sink_ready         (limiter_cmd_src_ready),             //       sink.ready
		.sink_channel       (limiter_cmd_src_channel),           //           .channel
		.sink_data          (limiter_cmd_src_data),              //           .data
		.sink_startofpacket (limiter_cmd_src_startofpacket),     //           .startofpacket
		.sink_endofpacket   (limiter_cmd_src_endofpacket),       //           .endofpacket
		.sink_valid         (limiter_cmd_valid_data),            // sink_valid.data
		.src0_ready         (cmd_xbar_demux_src0_ready),         //       src0.ready
		.src0_valid         (cmd_xbar_demux_src0_valid),         //           .valid
		.src0_data          (cmd_xbar_demux_src0_data),          //           .data
		.src0_channel       (cmd_xbar_demux_src0_channel),       //           .channel
		.src0_startofpacket (cmd_xbar_demux_src0_startofpacket), //           .startofpacket
		.src0_endofpacket   (cmd_xbar_demux_src0_endofpacket),   //           .endofpacket
		.src1_ready         (cmd_xbar_demux_src1_ready),         //       src1.ready
		.src1_valid         (cmd_xbar_demux_src1_valid),         //           .valid
		.src1_data          (cmd_xbar_demux_src1_data),          //           .data
		.src1_channel       (cmd_xbar_demux_src1_channel),       //           .channel
		.src1_startofpacket (cmd_xbar_demux_src1_startofpacket), //           .startofpacket
		.src1_endofpacket   (cmd_xbar_demux_src1_endofpacket)    //           .endofpacket
	);

	Nios1_cmd_xbar_demux_001 cmd_xbar_demux_001 (
		.clk                 (clk_clk),                                //        clk.clk
		.reset               (rst_controller_reset_out_reset),         //  clk_reset.reset
		.sink_ready          (limiter_001_cmd_src_ready),              //       sink.ready
		.sink_channel        (limiter_001_cmd_src_channel),            //           .channel
		.sink_data           (limiter_001_cmd_src_data),               //           .data
		.sink_startofpacket  (limiter_001_cmd_src_startofpacket),      //           .startofpacket
		.sink_endofpacket    (limiter_001_cmd_src_endofpacket),        //           .endofpacket
		.sink_valid          (limiter_001_cmd_valid_data),             // sink_valid.data
		.src0_ready          (cmd_xbar_demux_001_src0_ready),          //       src0.ready
		.src0_valid          (cmd_xbar_demux_001_src0_valid),          //           .valid
		.src0_data           (cmd_xbar_demux_001_src0_data),           //           .data
		.src0_channel        (cmd_xbar_demux_001_src0_channel),        //           .channel
		.src0_startofpacket  (cmd_xbar_demux_001_src0_startofpacket),  //           .startofpacket
		.src0_endofpacket    (cmd_xbar_demux_001_src0_endofpacket),    //           .endofpacket
		.src1_ready          (cmd_xbar_demux_001_src1_ready),          //       src1.ready
		.src1_valid          (cmd_xbar_demux_001_src1_valid),          //           .valid
		.src1_data           (cmd_xbar_demux_001_src1_data),           //           .data
		.src1_channel        (cmd_xbar_demux_001_src1_channel),        //           .channel
		.src1_startofpacket  (cmd_xbar_demux_001_src1_startofpacket),  //           .startofpacket
		.src1_endofpacket    (cmd_xbar_demux_001_src1_endofpacket),    //           .endofpacket
		.src2_ready          (cmd_xbar_demux_001_src2_ready),          //       src2.ready
		.src2_valid          (cmd_xbar_demux_001_src2_valid),          //           .valid
		.src2_data           (cmd_xbar_demux_001_src2_data),           //           .data
		.src2_channel        (cmd_xbar_demux_001_src2_channel),        //           .channel
		.src2_startofpacket  (cmd_xbar_demux_001_src2_startofpacket),  //           .startofpacket
		.src2_endofpacket    (cmd_xbar_demux_001_src2_endofpacket),    //           .endofpacket
		.src3_ready          (cmd_xbar_demux_001_src3_ready),          //       src3.ready
		.src3_valid          (cmd_xbar_demux_001_src3_valid),          //           .valid
		.src3_data           (cmd_xbar_demux_001_src3_data),           //           .data
		.src3_channel        (cmd_xbar_demux_001_src3_channel),        //           .channel
		.src3_startofpacket  (cmd_xbar_demux_001_src3_startofpacket),  //           .startofpacket
		.src3_endofpacket    (cmd_xbar_demux_001_src3_endofpacket),    //           .endofpacket
		.src4_ready          (cmd_xbar_demux_001_src4_ready),          //       src4.ready
		.src4_valid          (cmd_xbar_demux_001_src4_valid),          //           .valid
		.src4_data           (cmd_xbar_demux_001_src4_data),           //           .data
		.src4_channel        (cmd_xbar_demux_001_src4_channel),        //           .channel
		.src4_startofpacket  (cmd_xbar_demux_001_src4_startofpacket),  //           .startofpacket
		.src4_endofpacket    (cmd_xbar_demux_001_src4_endofpacket),    //           .endofpacket
		.src5_ready          (cmd_xbar_demux_001_src5_ready),          //       src5.ready
		.src5_valid          (cmd_xbar_demux_001_src5_valid),          //           .valid
		.src5_data           (cmd_xbar_demux_001_src5_data),           //           .data
		.src5_channel        (cmd_xbar_demux_001_src5_channel),        //           .channel
		.src5_startofpacket  (cmd_xbar_demux_001_src5_startofpacket),  //           .startofpacket
		.src5_endofpacket    (cmd_xbar_demux_001_src5_endofpacket),    //           .endofpacket
		.src6_ready          (cmd_xbar_demux_001_src6_ready),          //       src6.ready
		.src6_valid          (cmd_xbar_demux_001_src6_valid),          //           .valid
		.src6_data           (cmd_xbar_demux_001_src6_data),           //           .data
		.src6_channel        (cmd_xbar_demux_001_src6_channel),        //           .channel
		.src6_startofpacket  (cmd_xbar_demux_001_src6_startofpacket),  //           .startofpacket
		.src6_endofpacket    (cmd_xbar_demux_001_src6_endofpacket),    //           .endofpacket
		.src7_ready          (cmd_xbar_demux_001_src7_ready),          //       src7.ready
		.src7_valid          (cmd_xbar_demux_001_src7_valid),          //           .valid
		.src7_data           (cmd_xbar_demux_001_src7_data),           //           .data
		.src7_channel        (cmd_xbar_demux_001_src7_channel),        //           .channel
		.src7_startofpacket  (cmd_xbar_demux_001_src7_startofpacket),  //           .startofpacket
		.src7_endofpacket    (cmd_xbar_demux_001_src7_endofpacket),    //           .endofpacket
		.src8_ready          (cmd_xbar_demux_001_src8_ready),          //       src8.ready
		.src8_valid          (cmd_xbar_demux_001_src8_valid),          //           .valid
		.src8_data           (cmd_xbar_demux_001_src8_data),           //           .data
		.src8_channel        (cmd_xbar_demux_001_src8_channel),        //           .channel
		.src8_startofpacket  (cmd_xbar_demux_001_src8_startofpacket),  //           .startofpacket
		.src8_endofpacket    (cmd_xbar_demux_001_src8_endofpacket),    //           .endofpacket
		.src9_ready          (cmd_xbar_demux_001_src9_ready),          //       src9.ready
		.src9_valid          (cmd_xbar_demux_001_src9_valid),          //           .valid
		.src9_data           (cmd_xbar_demux_001_src9_data),           //           .data
		.src9_channel        (cmd_xbar_demux_001_src9_channel),        //           .channel
		.src9_startofpacket  (cmd_xbar_demux_001_src9_startofpacket),  //           .startofpacket
		.src9_endofpacket    (cmd_xbar_demux_001_src9_endofpacket),    //           .endofpacket
		.src10_ready         (cmd_xbar_demux_001_src10_ready),         //      src10.ready
		.src10_valid         (cmd_xbar_demux_001_src10_valid),         //           .valid
		.src10_data          (cmd_xbar_demux_001_src10_data),          //           .data
		.src10_channel       (cmd_xbar_demux_001_src10_channel),       //           .channel
		.src10_startofpacket (cmd_xbar_demux_001_src10_startofpacket), //           .startofpacket
		.src10_endofpacket   (cmd_xbar_demux_001_src10_endofpacket),   //           .endofpacket
		.src11_ready         (cmd_xbar_demux_001_src11_ready),         //      src11.ready
		.src11_valid         (cmd_xbar_demux_001_src11_valid),         //           .valid
		.src11_data          (cmd_xbar_demux_001_src11_data),          //           .data
		.src11_channel       (cmd_xbar_demux_001_src11_channel),       //           .channel
		.src11_startofpacket (cmd_xbar_demux_001_src11_startofpacket), //           .startofpacket
		.src11_endofpacket   (cmd_xbar_demux_001_src11_endofpacket),   //           .endofpacket
		.src12_ready         (cmd_xbar_demux_001_src12_ready),         //      src12.ready
		.src12_valid         (cmd_xbar_demux_001_src12_valid),         //           .valid
		.src12_data          (cmd_xbar_demux_001_src12_data),          //           .data
		.src12_channel       (cmd_xbar_demux_001_src12_channel),       //           .channel
		.src12_startofpacket (cmd_xbar_demux_001_src12_startofpacket), //           .startofpacket
		.src12_endofpacket   (cmd_xbar_demux_001_src12_endofpacket),   //           .endofpacket
		.src13_ready         (cmd_xbar_demux_001_src13_ready),         //      src13.ready
		.src13_valid         (cmd_xbar_demux_001_src13_valid),         //           .valid
		.src13_data          (cmd_xbar_demux_001_src13_data),          //           .data
		.src13_channel       (cmd_xbar_demux_001_src13_channel),       //           .channel
		.src13_startofpacket (cmd_xbar_demux_001_src13_startofpacket), //           .startofpacket
		.src13_endofpacket   (cmd_xbar_demux_001_src13_endofpacket)    //           .endofpacket
	);

	Nios1_cmd_xbar_mux cmd_xbar_mux (
		.clk                 (clk_clk),                               //       clk.clk
		.reset               (rst_controller_reset_out_reset),        // clk_reset.reset
		.src_ready           (cmd_xbar_mux_src_ready),                //       src.ready
		.src_valid           (cmd_xbar_mux_src_valid),                //          .valid
		.src_data            (cmd_xbar_mux_src_data),                 //          .data
		.src_channel         (cmd_xbar_mux_src_channel),              //          .channel
		.src_startofpacket   (cmd_xbar_mux_src_startofpacket),        //          .startofpacket
		.src_endofpacket     (cmd_xbar_mux_src_endofpacket),          //          .endofpacket
		.sink0_ready         (cmd_xbar_demux_src0_ready),             //     sink0.ready
		.sink0_valid         (cmd_xbar_demux_src0_valid),             //          .valid
		.sink0_channel       (cmd_xbar_demux_src0_channel),           //          .channel
		.sink0_data          (cmd_xbar_demux_src0_data),              //          .data
		.sink0_startofpacket (cmd_xbar_demux_src0_startofpacket),     //          .startofpacket
		.sink0_endofpacket   (cmd_xbar_demux_src0_endofpacket),       //          .endofpacket
		.sink1_ready         (cmd_xbar_demux_001_src0_ready),         //     sink1.ready
		.sink1_valid         (cmd_xbar_demux_001_src0_valid),         //          .valid
		.sink1_channel       (cmd_xbar_demux_001_src0_channel),       //          .channel
		.sink1_data          (cmd_xbar_demux_001_src0_data),          //          .data
		.sink1_startofpacket (cmd_xbar_demux_001_src0_startofpacket), //          .startofpacket
		.sink1_endofpacket   (cmd_xbar_demux_001_src0_endofpacket)    //          .endofpacket
	);

	Nios1_cmd_xbar_mux cmd_xbar_mux_001 (
		.clk                 (clk_clk),                               //       clk.clk
		.reset               (rst_controller_reset_out_reset),        // clk_reset.reset
		.src_ready           (cmd_xbar_mux_001_src_ready),            //       src.ready
		.src_valid           (cmd_xbar_mux_001_src_valid),            //          .valid
		.src_data            (cmd_xbar_mux_001_src_data),             //          .data
		.src_channel         (cmd_xbar_mux_001_src_channel),          //          .channel
		.src_startofpacket   (cmd_xbar_mux_001_src_startofpacket),    //          .startofpacket
		.src_endofpacket     (cmd_xbar_mux_001_src_endofpacket),      //          .endofpacket
		.sink0_ready         (cmd_xbar_demux_src1_ready),             //     sink0.ready
		.sink0_valid         (cmd_xbar_demux_src1_valid),             //          .valid
		.sink0_channel       (cmd_xbar_demux_src1_channel),           //          .channel
		.sink0_data          (cmd_xbar_demux_src1_data),              //          .data
		.sink0_startofpacket (cmd_xbar_demux_src1_startofpacket),     //          .startofpacket
		.sink0_endofpacket   (cmd_xbar_demux_src1_endofpacket),       //          .endofpacket
		.sink1_ready         (cmd_xbar_demux_001_src1_ready),         //     sink1.ready
		.sink1_valid         (cmd_xbar_demux_001_src1_valid),         //          .valid
		.sink1_channel       (cmd_xbar_demux_001_src1_channel),       //          .channel
		.sink1_data          (cmd_xbar_demux_001_src1_data),          //          .data
		.sink1_startofpacket (cmd_xbar_demux_001_src1_startofpacket), //          .startofpacket
		.sink1_endofpacket   (cmd_xbar_demux_001_src1_endofpacket)    //          .endofpacket
	);

	Nios1_rsp_xbar_demux rsp_xbar_demux (
		.clk                (clk_clk),                           //       clk.clk
		.reset              (rst_controller_reset_out_reset),    // clk_reset.reset
		.sink_ready         (id_router_src_ready),               //      sink.ready
		.sink_channel       (id_router_src_channel),             //          .channel
		.sink_data          (id_router_src_data),                //          .data
		.sink_startofpacket (id_router_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_src0_endofpacket),   //          .endofpacket
		.src1_ready         (rsp_xbar_demux_src1_ready),         //      src1.ready
		.src1_valid         (rsp_xbar_demux_src1_valid),         //          .valid
		.src1_data          (rsp_xbar_demux_src1_data),          //          .data
		.src1_channel       (rsp_xbar_demux_src1_channel),       //          .channel
		.src1_startofpacket (rsp_xbar_demux_src1_startofpacket), //          .startofpacket
		.src1_endofpacket   (rsp_xbar_demux_src1_endofpacket)    //          .endofpacket
	);

	Nios1_rsp_xbar_demux rsp_xbar_demux_001 (
		.clk                (clk_clk),                               //       clk.clk
		.reset              (rst_controller_reset_out_reset),        // clk_reset.reset
		.sink_ready         (id_router_001_src_ready),               //      sink.ready
		.sink_channel       (id_router_001_src_channel),             //          .channel
		.sink_data          (id_router_001_src_data),                //          .data
		.sink_startofpacket (id_router_001_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_001_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_001_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_001_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_001_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_001_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_001_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_001_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_001_src0_endofpacket),   //          .endofpacket
		.src1_ready         (rsp_xbar_demux_001_src1_ready),         //      src1.ready
		.src1_valid         (rsp_xbar_demux_001_src1_valid),         //          .valid
		.src1_data          (rsp_xbar_demux_001_src1_data),          //          .data
		.src1_channel       (rsp_xbar_demux_001_src1_channel),       //          .channel
		.src1_startofpacket (rsp_xbar_demux_001_src1_startofpacket), //          .startofpacket
		.src1_endofpacket   (rsp_xbar_demux_001_src1_endofpacket)    //          .endofpacket
	);

	Nios1_rsp_xbar_demux_002 rsp_xbar_demux_002 (
		.clk                (clk_clk),                               //       clk.clk
		.reset              (rst_controller_reset_out_reset),        // clk_reset.reset
		.sink_ready         (id_router_002_src_ready),               //      sink.ready
		.sink_channel       (id_router_002_src_channel),             //          .channel
		.sink_data          (id_router_002_src_data),                //          .data
		.sink_startofpacket (id_router_002_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_002_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_002_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_002_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_002_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_002_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_002_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_002_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_002_src0_endofpacket)    //          .endofpacket
	);

	Nios1_rsp_xbar_demux_002 rsp_xbar_demux_003 (
		.clk                (clk_clk),                               //       clk.clk
		.reset              (rst_controller_reset_out_reset),        // clk_reset.reset
		.sink_ready         (id_router_003_src_ready),               //      sink.ready
		.sink_channel       (id_router_003_src_channel),             //          .channel
		.sink_data          (id_router_003_src_data),                //          .data
		.sink_startofpacket (id_router_003_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_003_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_003_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_003_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_003_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_003_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_003_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_003_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_003_src0_endofpacket)    //          .endofpacket
	);

	Nios1_rsp_xbar_demux_002 rsp_xbar_demux_004 (
		.clk                (clk_clk),                               //       clk.clk
		.reset              (rst_controller_reset_out_reset),        // clk_reset.reset
		.sink_ready         (id_router_004_src_ready),               //      sink.ready
		.sink_channel       (id_router_004_src_channel),             //          .channel
		.sink_data          (id_router_004_src_data),                //          .data
		.sink_startofpacket (id_router_004_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_004_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_004_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_004_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_004_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_004_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_004_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_004_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_004_src0_endofpacket)    //          .endofpacket
	);

	Nios1_rsp_xbar_demux_002 rsp_xbar_demux_005 (
		.clk                (clk_clk),                               //       clk.clk
		.reset              (rst_controller_reset_out_reset),        // clk_reset.reset
		.sink_ready         (id_router_005_src_ready),               //      sink.ready
		.sink_channel       (id_router_005_src_channel),             //          .channel
		.sink_data          (id_router_005_src_data),                //          .data
		.sink_startofpacket (id_router_005_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_005_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_005_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_005_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_005_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_005_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_005_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_005_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_005_src0_endofpacket)    //          .endofpacket
	);

	Nios1_rsp_xbar_demux_002 rsp_xbar_demux_006 (
		.clk                (clk_clk),                               //       clk.clk
		.reset              (rst_controller_reset_out_reset),        // clk_reset.reset
		.sink_ready         (id_router_006_src_ready),               //      sink.ready
		.sink_channel       (id_router_006_src_channel),             //          .channel
		.sink_data          (id_router_006_src_data),                //          .data
		.sink_startofpacket (id_router_006_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_006_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_006_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_006_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_006_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_006_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_006_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_006_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_006_src0_endofpacket)    //          .endofpacket
	);

	Nios1_rsp_xbar_demux_002 rsp_xbar_demux_007 (
		.clk                (clk_clk),                               //       clk.clk
		.reset              (rst_controller_reset_out_reset),        // clk_reset.reset
		.sink_ready         (id_router_007_src_ready),               //      sink.ready
		.sink_channel       (id_router_007_src_channel),             //          .channel
		.sink_data          (id_router_007_src_data),                //          .data
		.sink_startofpacket (id_router_007_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_007_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_007_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_007_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_007_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_007_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_007_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_007_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_007_src0_endofpacket)    //          .endofpacket
	);

	Nios1_rsp_xbar_demux_002 rsp_xbar_demux_008 (
		.clk                (clk_clk),                               //       clk.clk
		.reset              (rst_controller_reset_out_reset),        // clk_reset.reset
		.sink_ready         (id_router_008_src_ready),               //      sink.ready
		.sink_channel       (id_router_008_src_channel),             //          .channel
		.sink_data          (id_router_008_src_data),                //          .data
		.sink_startofpacket (id_router_008_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_008_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_008_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_008_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_008_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_008_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_008_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_008_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_008_src0_endofpacket)    //          .endofpacket
	);

	Nios1_rsp_xbar_demux_002 rsp_xbar_demux_009 (
		.clk                (clk_clk),                               //       clk.clk
		.reset              (rst_controller_reset_out_reset),        // clk_reset.reset
		.sink_ready         (id_router_009_src_ready),               //      sink.ready
		.sink_channel       (id_router_009_src_channel),             //          .channel
		.sink_data          (id_router_009_src_data),                //          .data
		.sink_startofpacket (id_router_009_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_009_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_009_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_009_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_009_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_009_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_009_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_009_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_009_src0_endofpacket)    //          .endofpacket
	);

	Nios1_rsp_xbar_demux_002 rsp_xbar_demux_010 (
		.clk                (clk_clk),                               //       clk.clk
		.reset              (rst_controller_reset_out_reset),        // clk_reset.reset
		.sink_ready         (id_router_010_src_ready),               //      sink.ready
		.sink_channel       (id_router_010_src_channel),             //          .channel
		.sink_data          (id_router_010_src_data),                //          .data
		.sink_startofpacket (id_router_010_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_010_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_010_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_010_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_010_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_010_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_010_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_010_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_010_src0_endofpacket)    //          .endofpacket
	);

	Nios1_rsp_xbar_demux_002 rsp_xbar_demux_011 (
		.clk                (clk_clk),                               //       clk.clk
		.reset              (rst_controller_reset_out_reset),        // clk_reset.reset
		.sink_ready         (id_router_011_src_ready),               //      sink.ready
		.sink_channel       (id_router_011_src_channel),             //          .channel
		.sink_data          (id_router_011_src_data),                //          .data
		.sink_startofpacket (id_router_011_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_011_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_011_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_011_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_011_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_011_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_011_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_011_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_011_src0_endofpacket)    //          .endofpacket
	);

	Nios1_rsp_xbar_demux_002 rsp_xbar_demux_012 (
		.clk                (clk_clk),                               //       clk.clk
		.reset              (rst_controller_reset_out_reset),        // clk_reset.reset
		.sink_ready         (id_router_012_src_ready),               //      sink.ready
		.sink_channel       (id_router_012_src_channel),             //          .channel
		.sink_data          (id_router_012_src_data),                //          .data
		.sink_startofpacket (id_router_012_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_012_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_012_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_012_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_012_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_012_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_012_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_012_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_012_src0_endofpacket)    //          .endofpacket
	);

	Nios1_rsp_xbar_demux_002 rsp_xbar_demux_013 (
		.clk                (clk_clk),                               //       clk.clk
		.reset              (rst_controller_reset_out_reset),        // clk_reset.reset
		.sink_ready         (id_router_013_src_ready),               //      sink.ready
		.sink_channel       (id_router_013_src_channel),             //          .channel
		.sink_data          (id_router_013_src_data),                //          .data
		.sink_startofpacket (id_router_013_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_013_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_013_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_013_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_013_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_013_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_013_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_013_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_013_src0_endofpacket)    //          .endofpacket
	);

	Nios1_rsp_xbar_mux rsp_xbar_mux (
		.clk                 (clk_clk),                               //       clk.clk
		.reset               (rst_controller_reset_out_reset),        // clk_reset.reset
		.src_ready           (rsp_xbar_mux_src_ready),                //       src.ready
		.src_valid           (rsp_xbar_mux_src_valid),                //          .valid
		.src_data            (rsp_xbar_mux_src_data),                 //          .data
		.src_channel         (rsp_xbar_mux_src_channel),              //          .channel
		.src_startofpacket   (rsp_xbar_mux_src_startofpacket),        //          .startofpacket
		.src_endofpacket     (rsp_xbar_mux_src_endofpacket),          //          .endofpacket
		.sink0_ready         (rsp_xbar_demux_src0_ready),             //     sink0.ready
		.sink0_valid         (rsp_xbar_demux_src0_valid),             //          .valid
		.sink0_channel       (rsp_xbar_demux_src0_channel),           //          .channel
		.sink0_data          (rsp_xbar_demux_src0_data),              //          .data
		.sink0_startofpacket (rsp_xbar_demux_src0_startofpacket),     //          .startofpacket
		.sink0_endofpacket   (rsp_xbar_demux_src0_endofpacket),       //          .endofpacket
		.sink1_ready         (rsp_xbar_demux_001_src0_ready),         //     sink1.ready
		.sink1_valid         (rsp_xbar_demux_001_src0_valid),         //          .valid
		.sink1_channel       (rsp_xbar_demux_001_src0_channel),       //          .channel
		.sink1_data          (rsp_xbar_demux_001_src0_data),          //          .data
		.sink1_startofpacket (rsp_xbar_demux_001_src0_startofpacket), //          .startofpacket
		.sink1_endofpacket   (rsp_xbar_demux_001_src0_endofpacket)    //          .endofpacket
	);

	Nios1_rsp_xbar_mux_001 rsp_xbar_mux_001 (
		.clk                  (clk_clk),                               //       clk.clk
		.reset                (rst_controller_reset_out_reset),        // clk_reset.reset
		.src_ready            (rsp_xbar_mux_001_src_ready),            //       src.ready
		.src_valid            (rsp_xbar_mux_001_src_valid),            //          .valid
		.src_data             (rsp_xbar_mux_001_src_data),             //          .data
		.src_channel          (rsp_xbar_mux_001_src_channel),          //          .channel
		.src_startofpacket    (rsp_xbar_mux_001_src_startofpacket),    //          .startofpacket
		.src_endofpacket      (rsp_xbar_mux_001_src_endofpacket),      //          .endofpacket
		.sink0_ready          (rsp_xbar_demux_src1_ready),             //     sink0.ready
		.sink0_valid          (rsp_xbar_demux_src1_valid),             //          .valid
		.sink0_channel        (rsp_xbar_demux_src1_channel),           //          .channel
		.sink0_data           (rsp_xbar_demux_src1_data),              //          .data
		.sink0_startofpacket  (rsp_xbar_demux_src1_startofpacket),     //          .startofpacket
		.sink0_endofpacket    (rsp_xbar_demux_src1_endofpacket),       //          .endofpacket
		.sink1_ready          (rsp_xbar_demux_001_src1_ready),         //     sink1.ready
		.sink1_valid          (rsp_xbar_demux_001_src1_valid),         //          .valid
		.sink1_channel        (rsp_xbar_demux_001_src1_channel),       //          .channel
		.sink1_data           (rsp_xbar_demux_001_src1_data),          //          .data
		.sink1_startofpacket  (rsp_xbar_demux_001_src1_startofpacket), //          .startofpacket
		.sink1_endofpacket    (rsp_xbar_demux_001_src1_endofpacket),   //          .endofpacket
		.sink2_ready          (rsp_xbar_demux_002_src0_ready),         //     sink2.ready
		.sink2_valid          (rsp_xbar_demux_002_src0_valid),         //          .valid
		.sink2_channel        (rsp_xbar_demux_002_src0_channel),       //          .channel
		.sink2_data           (rsp_xbar_demux_002_src0_data),          //          .data
		.sink2_startofpacket  (rsp_xbar_demux_002_src0_startofpacket), //          .startofpacket
		.sink2_endofpacket    (rsp_xbar_demux_002_src0_endofpacket),   //          .endofpacket
		.sink3_ready          (rsp_xbar_demux_003_src0_ready),         //     sink3.ready
		.sink3_valid          (rsp_xbar_demux_003_src0_valid),         //          .valid
		.sink3_channel        (rsp_xbar_demux_003_src0_channel),       //          .channel
		.sink3_data           (rsp_xbar_demux_003_src0_data),          //          .data
		.sink3_startofpacket  (rsp_xbar_demux_003_src0_startofpacket), //          .startofpacket
		.sink3_endofpacket    (rsp_xbar_demux_003_src0_endofpacket),   //          .endofpacket
		.sink4_ready          (rsp_xbar_demux_004_src0_ready),         //     sink4.ready
		.sink4_valid          (rsp_xbar_demux_004_src0_valid),         //          .valid
		.sink4_channel        (rsp_xbar_demux_004_src0_channel),       //          .channel
		.sink4_data           (rsp_xbar_demux_004_src0_data),          //          .data
		.sink4_startofpacket  (rsp_xbar_demux_004_src0_startofpacket), //          .startofpacket
		.sink4_endofpacket    (rsp_xbar_demux_004_src0_endofpacket),   //          .endofpacket
		.sink5_ready          (rsp_xbar_demux_005_src0_ready),         //     sink5.ready
		.sink5_valid          (rsp_xbar_demux_005_src0_valid),         //          .valid
		.sink5_channel        (rsp_xbar_demux_005_src0_channel),       //          .channel
		.sink5_data           (rsp_xbar_demux_005_src0_data),          //          .data
		.sink5_startofpacket  (rsp_xbar_demux_005_src0_startofpacket), //          .startofpacket
		.sink5_endofpacket    (rsp_xbar_demux_005_src0_endofpacket),   //          .endofpacket
		.sink6_ready          (rsp_xbar_demux_006_src0_ready),         //     sink6.ready
		.sink6_valid          (rsp_xbar_demux_006_src0_valid),         //          .valid
		.sink6_channel        (rsp_xbar_demux_006_src0_channel),       //          .channel
		.sink6_data           (rsp_xbar_demux_006_src0_data),          //          .data
		.sink6_startofpacket  (rsp_xbar_demux_006_src0_startofpacket), //          .startofpacket
		.sink6_endofpacket    (rsp_xbar_demux_006_src0_endofpacket),   //          .endofpacket
		.sink7_ready          (rsp_xbar_demux_007_src0_ready),         //     sink7.ready
		.sink7_valid          (rsp_xbar_demux_007_src0_valid),         //          .valid
		.sink7_channel        (rsp_xbar_demux_007_src0_channel),       //          .channel
		.sink7_data           (rsp_xbar_demux_007_src0_data),          //          .data
		.sink7_startofpacket  (rsp_xbar_demux_007_src0_startofpacket), //          .startofpacket
		.sink7_endofpacket    (rsp_xbar_demux_007_src0_endofpacket),   //          .endofpacket
		.sink8_ready          (rsp_xbar_demux_008_src0_ready),         //     sink8.ready
		.sink8_valid          (rsp_xbar_demux_008_src0_valid),         //          .valid
		.sink8_channel        (rsp_xbar_demux_008_src0_channel),       //          .channel
		.sink8_data           (rsp_xbar_demux_008_src0_data),          //          .data
		.sink8_startofpacket  (rsp_xbar_demux_008_src0_startofpacket), //          .startofpacket
		.sink8_endofpacket    (rsp_xbar_demux_008_src0_endofpacket),   //          .endofpacket
		.sink9_ready          (rsp_xbar_demux_009_src0_ready),         //     sink9.ready
		.sink9_valid          (rsp_xbar_demux_009_src0_valid),         //          .valid
		.sink9_channel        (rsp_xbar_demux_009_src0_channel),       //          .channel
		.sink9_data           (rsp_xbar_demux_009_src0_data),          //          .data
		.sink9_startofpacket  (rsp_xbar_demux_009_src0_startofpacket), //          .startofpacket
		.sink9_endofpacket    (rsp_xbar_demux_009_src0_endofpacket),   //          .endofpacket
		.sink10_ready         (rsp_xbar_demux_010_src0_ready),         //    sink10.ready
		.sink10_valid         (rsp_xbar_demux_010_src0_valid),         //          .valid
		.sink10_channel       (rsp_xbar_demux_010_src0_channel),       //          .channel
		.sink10_data          (rsp_xbar_demux_010_src0_data),          //          .data
		.sink10_startofpacket (rsp_xbar_demux_010_src0_startofpacket), //          .startofpacket
		.sink10_endofpacket   (rsp_xbar_demux_010_src0_endofpacket),   //          .endofpacket
		.sink11_ready         (rsp_xbar_demux_011_src0_ready),         //    sink11.ready
		.sink11_valid         (rsp_xbar_demux_011_src0_valid),         //          .valid
		.sink11_channel       (rsp_xbar_demux_011_src0_channel),       //          .channel
		.sink11_data          (rsp_xbar_demux_011_src0_data),          //          .data
		.sink11_startofpacket (rsp_xbar_demux_011_src0_startofpacket), //          .startofpacket
		.sink11_endofpacket   (rsp_xbar_demux_011_src0_endofpacket),   //          .endofpacket
		.sink12_ready         (rsp_xbar_demux_012_src0_ready),         //    sink12.ready
		.sink12_valid         (rsp_xbar_demux_012_src0_valid),         //          .valid
		.sink12_channel       (rsp_xbar_demux_012_src0_channel),       //          .channel
		.sink12_data          (rsp_xbar_demux_012_src0_data),          //          .data
		.sink12_startofpacket (rsp_xbar_demux_012_src0_startofpacket), //          .startofpacket
		.sink12_endofpacket   (rsp_xbar_demux_012_src0_endofpacket),   //          .endofpacket
		.sink13_ready         (rsp_xbar_demux_013_src0_ready),         //    sink13.ready
		.sink13_valid         (rsp_xbar_demux_013_src0_valid),         //          .valid
		.sink13_channel       (rsp_xbar_demux_013_src0_channel),       //          .channel
		.sink13_data          (rsp_xbar_demux_013_src0_data),          //          .data
		.sink13_startofpacket (rsp_xbar_demux_013_src0_startofpacket), //          .startofpacket
		.sink13_endofpacket   (rsp_xbar_demux_013_src0_endofpacket)    //          .endofpacket
	);

	Nios1_irq_mapper irq_mapper (
		.clk           (clk_clk),                        //       clk.clk
		.reset         (rst_controller_reset_out_reset), // clk_reset.reset
		.receiver0_irq (irq_mapper_receiver0_irq),       // receiver0.irq
		.receiver1_irq (irq_mapper_receiver1_irq),       // receiver1.irq
		.receiver2_irq (irq_mapper_receiver2_irq),       // receiver2.irq
		.receiver3_irq (irq_mapper_receiver3_irq),       // receiver3.irq
		.receiver4_irq (irq_mapper_receiver4_irq),       // receiver4.irq
		.sender_irq    (nios2_qsys_d_irq_irq)            //    sender.irq
	);

endmodule
