-- Nios1.vhd

-- Generated using ACDS version 11.1sp2 259 at 2012.10.25.17:22:09

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity Nios1 is
	port (
		pio_ledr_export     : out   std_logic_vector(17 downto 0);                    --      pio_ledr.export
		pio_dataread_export : out   std_logic_vector(1 downto 0);                     --  pio_dataread.export
		pio_data_export     : in    std_logic_vector(11 downto 0) := (others => '0'); --      pio_data.export
		pio_ledg_export     : out   std_logic_vector(7 downto 0);                     --      pio_ledg.export
		pio_sw_export       : in    std_logic_vector(17 downto 0) := (others => '0'); --        pio_sw.export
		uart_external_rxd   : in    std_logic                     := '0';             -- uart_external.rxd
		uart_external_txd   : out   std_logic;                                        --              .txd
		pio_rdydata_export  : in    std_logic                     := '0';             --   pio_rdydata.export
		lcd_external_data   : inout std_logic_vector(7 downto 0)  := (others => '0'); --  lcd_external.data
		lcd_external_E      : out   std_logic;                                        --              .E
		lcd_external_RS     : out   std_logic;                                        --              .RS
		lcd_external_RW     : out   std_logic;                                        --              .RW
		reset_reset_n       : in    std_logic                     := '0';             --         reset.reset_n
		clk_clk             : in    std_logic                     := '0';             --           clk.clk
		pio_button_export   : in    std_logic_vector(2 downto 0)  := (others => '0')  --    pio_button.export
	);
end entity Nios1;

architecture rtl of Nios1 is
	component Nios1_nios2_qsys is
		port (
			clk                                   : in  std_logic                     := 'X';             -- clk
			reset_n                               : in  std_logic                     := 'X';             -- reset_n
			d_address                             : out std_logic_vector(18 downto 0);                    -- address
			d_byteenable                          : out std_logic_vector(3 downto 0);                     -- byteenable
			d_read                                : out std_logic;                                        -- read
			d_readdata                            : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			d_waitrequest                         : in  std_logic                     := 'X';             -- waitrequest
			d_write                               : out std_logic;                                        -- write
			d_writedata                           : out std_logic_vector(31 downto 0);                    -- writedata
			d_readdatavalid                       : in  std_logic                     := 'X';             -- readdatavalid
			jtag_debug_module_debugaccess_to_roms : out std_logic;                                        -- debugaccess
			i_address                             : out std_logic_vector(18 downto 0);                    -- address
			i_read                                : out std_logic;                                        -- read
			i_readdata                            : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			i_waitrequest                         : in  std_logic                     := 'X';             -- waitrequest
			i_readdatavalid                       : in  std_logic                     := 'X';             -- readdatavalid
			d_irq                                 : in  std_logic_vector(31 downto 0) := (others => 'X'); -- irq
			jtag_debug_module_resetrequest        : out std_logic;                                        -- reset
			jtag_debug_module_address             : in  std_logic_vector(8 downto 0)  := (others => 'X'); -- address
			jtag_debug_module_begintransfer       : in  std_logic                     := 'X';             -- begintransfer
			jtag_debug_module_byteenable          : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			jtag_debug_module_debugaccess         : in  std_logic                     := 'X';             -- debugaccess
			jtag_debug_module_readdata            : out std_logic_vector(31 downto 0);                    -- readdata
			jtag_debug_module_select              : in  std_logic                     := 'X';             -- chipselect
			jtag_debug_module_write               : in  std_logic                     := 'X';             -- write
			jtag_debug_module_writedata           : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			no_ci_readra                          : out std_logic                                         -- readra
		);
	end component Nios1_nios2_qsys;

	component Nios1_onchip_memory is
		port (
			clk        : in  std_logic                     := 'X';             -- clk
			address    : in  std_logic_vector(14 downto 0) := (others => 'X'); -- address
			chipselect : in  std_logic                     := 'X';             -- chipselect
			clken      : in  std_logic                     := 'X';             -- clken
			readdata   : out std_logic_vector(31 downto 0);                    -- readdata
			write      : in  std_logic                     := 'X';             -- write
			writedata  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			byteenable : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			reset      : in  std_logic                     := 'X'              -- reset
		);
	end component Nios1_onchip_memory;

	component Nios1_jtag_uart is
		port (
			clk            : in  std_logic                     := 'X';             -- clk
			rst_n          : in  std_logic                     := 'X';             -- reset_n
			av_chipselect  : in  std_logic                     := 'X';             -- chipselect
			av_address     : in  std_logic                     := 'X';             -- address
			av_read_n      : in  std_logic                     := 'X';             -- read_n
			av_readdata    : out std_logic_vector(31 downto 0);                    -- readdata
			av_write_n     : in  std_logic                     := 'X';             -- write_n
			av_writedata   : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			av_waitrequest : out std_logic;                                        -- waitrequest
			dataavailable  : out std_logic;                                        -- dataavailable
			readyfordata   : out std_logic;                                        -- readyfordata
			av_irq         : out std_logic                                         -- irq
		);
	end component Nios1_jtag_uart;

	component Nios1_sysid_qsys is
		port (
			clock    : in  std_logic                     := 'X'; -- clk
			reset_n  : in  std_logic                     := 'X'; -- reset_n
			readdata : out std_logic_vector(31 downto 0);        -- readdata
			address  : in  std_logic                     := 'X'  -- address
		);
	end component Nios1_sysid_qsys;

	component Nios1_pio_LEDG is
		port (
			clk        : in  std_logic                     := 'X';             -- clk
			reset_n    : in  std_logic                     := 'X';             -- reset_n
			address    : in  std_logic_vector(2 downto 0)  := (others => 'X'); -- address
			write_n    : in  std_logic                     := 'X';             -- write_n
			writedata  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			chipselect : in  std_logic                     := 'X';             -- chipselect
			readdata   : out std_logic_vector(31 downto 0);                    -- readdata
			out_port   : out std_logic_vector(7 downto 0)                      -- export
		);
	end component Nios1_pio_LEDG;

	component Nios1_pio_LEDR is
		port (
			clk        : in  std_logic                     := 'X';             -- clk
			reset_n    : in  std_logic                     := 'X';             -- reset_n
			address    : in  std_logic_vector(2 downto 0)  := (others => 'X'); -- address
			write_n    : in  std_logic                     := 'X';             -- write_n
			writedata  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			chipselect : in  std_logic                     := 'X';             -- chipselect
			readdata   : out std_logic_vector(31 downto 0);                    -- readdata
			out_port   : out std_logic_vector(17 downto 0)                     -- export
		);
	end component Nios1_pio_LEDR;

	component Nios1_pio_SW is
		port (
			clk      : in  std_logic                     := 'X';             -- clk
			reset_n  : in  std_logic                     := 'X';             -- reset_n
			address  : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- address
			readdata : out std_logic_vector(31 downto 0);                    -- readdata
			in_port  : in  std_logic_vector(17 downto 0) := (others => 'X')  -- export
		);
	end component Nios1_pio_SW;

	component Nios1_pio_Button is
		port (
			clk        : in  std_logic                     := 'X';             -- clk
			reset_n    : in  std_logic                     := 'X';             -- reset_n
			address    : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- address
			write_n    : in  std_logic                     := 'X';             -- write_n
			writedata  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			chipselect : in  std_logic                     := 'X';             -- chipselect
			readdata   : out std_logic_vector(31 downto 0);                    -- readdata
			in_port    : in  std_logic_vector(2 downto 0)  := (others => 'X'); -- export
			irq        : out std_logic                                         -- irq
		);
	end component Nios1_pio_Button;

	component Nios1_lcd is
		port (
			clk           : in    std_logic                    := 'X';             -- clk
			reset_n       : in    std_logic                    := 'X';             -- reset_n
			address       : in    std_logic_vector(1 downto 0) := (others => 'X'); -- address
			begintransfer : in    std_logic                    := 'X';             -- begintransfer
			read          : in    std_logic                    := 'X';             -- read
			readdata      : out   std_logic_vector(7 downto 0);                    -- readdata
			write         : in    std_logic                    := 'X';             -- write
			writedata     : in    std_logic_vector(7 downto 0) := (others => 'X'); -- writedata
			LCD_data      : inout std_logic_vector(7 downto 0) := (others => 'X'); -- export
			LCD_E         : out   std_logic;                                       -- export
			LCD_RS        : out   std_logic;                                       -- export
			LCD_RW        : out   std_logic                                        -- export
		);
	end component Nios1_lcd;

	component Nios1_uart is
		port (
			clk           : in  std_logic                     := 'X';             -- clk
			reset_n       : in  std_logic                     := 'X';             -- reset_n
			address       : in  std_logic_vector(2 downto 0)  := (others => 'X'); -- address
			begintransfer : in  std_logic                     := 'X';             -- begintransfer
			chipselect    : in  std_logic                     := 'X';             -- chipselect
			read_n        : in  std_logic                     := 'X';             -- read_n
			write_n       : in  std_logic                     := 'X';             -- write_n
			writedata     : in  std_logic_vector(15 downto 0) := (others => 'X'); -- writedata
			readdata      : out std_logic_vector(15 downto 0);                    -- readdata
			dataavailable : out std_logic;                                        -- dataavailable
			readyfordata  : out std_logic;                                        -- readyfordata
			rxd           : in  std_logic                     := 'X';             -- export
			txd           : out std_logic;                                        -- export
			irq           : out std_logic                                         -- irq
		);
	end component Nios1_uart;

	component Nios1_timer_0 is
		port (
			clk        : in  std_logic                     := 'X';             -- clk
			reset_n    : in  std_logic                     := 'X';             -- reset_n
			address    : in  std_logic_vector(2 downto 0)  := (others => 'X'); -- address
			writedata  : in  std_logic_vector(15 downto 0) := (others => 'X'); -- writedata
			readdata   : out std_logic_vector(15 downto 0);                    -- readdata
			chipselect : in  std_logic                     := 'X';             -- chipselect
			write_n    : in  std_logic                     := 'X';             -- write_n
			irq        : out std_logic                                         -- irq
		);
	end component Nios1_timer_0;

	component Nios1_pio_Data is
		port (
			clk      : in  std_logic                     := 'X';             -- clk
			reset_n  : in  std_logic                     := 'X';             -- reset_n
			address  : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- address
			readdata : out std_logic_vector(31 downto 0);                    -- readdata
			in_port  : in  std_logic_vector(11 downto 0) := (others => 'X')  -- export
		);
	end component Nios1_pio_Data;

	component Nios1_pio_RdyData is
		port (
			clk        : in  std_logic                     := 'X';             -- clk
			reset_n    : in  std_logic                     := 'X';             -- reset_n
			address    : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- address
			write_n    : in  std_logic                     := 'X';             -- write_n
			writedata  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			chipselect : in  std_logic                     := 'X';             -- chipselect
			readdata   : out std_logic_vector(31 downto 0);                    -- readdata
			in_port    : in  std_logic                     := 'X';             -- export
			irq        : out std_logic                                         -- irq
		);
	end component Nios1_pio_RdyData;

	component Nios1_pio_DataRead is
		port (
			clk        : in  std_logic                     := 'X';             -- clk
			reset_n    : in  std_logic                     := 'X';             -- reset_n
			address    : in  std_logic_vector(2 downto 0)  := (others => 'X'); -- address
			write_n    : in  std_logic                     := 'X';             -- write_n
			writedata  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			chipselect : in  std_logic                     := 'X';             -- chipselect
			readdata   : out std_logic_vector(31 downto 0);                    -- readdata
			out_port   : out std_logic_vector(1 downto 0)                      -- export
		);
	end component Nios1_pio_DataRead;

	component Nios1_nios2_qsys_instruction_master_translator is
		port (
			clk               : in  std_logic                     := 'X';             -- clk
			reset             : in  std_logic                     := 'X';             -- reset
			uav_address       : out std_logic_vector(18 downto 0);                    -- address
			uav_burstcount    : out std_logic_vector(2 downto 0);                     -- burstcount
			uav_read          : out std_logic;                                        -- read
			uav_write         : out std_logic;                                        -- write
			uav_waitrequest   : in  std_logic                     := 'X';             -- waitrequest
			uav_readdatavalid : in  std_logic                     := 'X';             -- readdatavalid
			uav_byteenable    : out std_logic_vector(3 downto 0);                     -- byteenable
			uav_readdata      : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			uav_writedata     : out std_logic_vector(31 downto 0);                    -- writedata
			uav_lock          : out std_logic;                                        -- lock
			uav_debugaccess   : out std_logic;                                        -- debugaccess
			av_address        : in  std_logic_vector(18 downto 0) := (others => 'X'); -- address
			av_waitrequest    : out std_logic;                                        -- waitrequest
			av_read           : in  std_logic                     := 'X';             -- read
			av_readdata       : out std_logic_vector(31 downto 0);                    -- readdata
			av_readdatavalid  : out std_logic                                         -- readdatavalid
		);
	end component Nios1_nios2_qsys_instruction_master_translator;

	component Nios1_nios2_qsys_data_master_translator is
		port (
			clk               : in  std_logic                     := 'X';             -- clk
			reset             : in  std_logic                     := 'X';             -- reset
			uav_address       : out std_logic_vector(18 downto 0);                    -- address
			uav_burstcount    : out std_logic_vector(2 downto 0);                     -- burstcount
			uav_read          : out std_logic;                                        -- read
			uav_write         : out std_logic;                                        -- write
			uav_waitrequest   : in  std_logic                     := 'X';             -- waitrequest
			uav_readdatavalid : in  std_logic                     := 'X';             -- readdatavalid
			uav_byteenable    : out std_logic_vector(3 downto 0);                     -- byteenable
			uav_readdata      : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			uav_writedata     : out std_logic_vector(31 downto 0);                    -- writedata
			uav_lock          : out std_logic;                                        -- lock
			uav_debugaccess   : out std_logic;                                        -- debugaccess
			av_address        : in  std_logic_vector(18 downto 0) := (others => 'X'); -- address
			av_waitrequest    : out std_logic;                                        -- waitrequest
			av_byteenable     : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			av_read           : in  std_logic                     := 'X';             -- read
			av_readdata       : out std_logic_vector(31 downto 0);                    -- readdata
			av_readdatavalid  : out std_logic;                                        -- readdatavalid
			av_write          : in  std_logic                     := 'X';             -- write
			av_writedata      : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			av_debugaccess    : in  std_logic                     := 'X'              -- debugaccess
		);
	end component Nios1_nios2_qsys_data_master_translator;

	component Nios1_nios2_qsys_jtag_debug_module_translator is
		port (
			clk               : in  std_logic                     := 'X';             -- clk
			reset             : in  std_logic                     := 'X';             -- reset
			uav_address       : in  std_logic_vector(18 downto 0) := (others => 'X'); -- address
			uav_burstcount    : in  std_logic_vector(2 downto 0)  := (others => 'X'); -- burstcount
			uav_read          : in  std_logic                     := 'X';             -- read
			uav_write         : in  std_logic                     := 'X';             -- write
			uav_waitrequest   : out std_logic;                                        -- waitrequest
			uav_readdatavalid : out std_logic;                                        -- readdatavalid
			uav_byteenable    : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			uav_readdata      : out std_logic_vector(31 downto 0);                    -- readdata
			uav_writedata     : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			uav_lock          : in  std_logic                     := 'X';             -- lock
			uav_debugaccess   : in  std_logic                     := 'X';             -- debugaccess
			av_address        : out std_logic_vector(8 downto 0);                     -- address
			av_write          : out std_logic;                                        -- write
			av_readdata       : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			av_writedata      : out std_logic_vector(31 downto 0);                    -- writedata
			av_begintransfer  : out std_logic;                                        -- begintransfer
			av_byteenable     : out std_logic_vector(3 downto 0);                     -- byteenable
			av_chipselect     : out std_logic;                                        -- chipselect
			av_debugaccess    : out std_logic                                         -- debugaccess
		);
	end component Nios1_nios2_qsys_jtag_debug_module_translator;

	component Nios1_onchip_memory_s1_translator is
		port (
			clk               : in  std_logic                     := 'X';             -- clk
			reset             : in  std_logic                     := 'X';             -- reset
			uav_address       : in  std_logic_vector(18 downto 0) := (others => 'X'); -- address
			uav_burstcount    : in  std_logic_vector(2 downto 0)  := (others => 'X'); -- burstcount
			uav_read          : in  std_logic                     := 'X';             -- read
			uav_write         : in  std_logic                     := 'X';             -- write
			uav_waitrequest   : out std_logic;                                        -- waitrequest
			uav_readdatavalid : out std_logic;                                        -- readdatavalid
			uav_byteenable    : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			uav_readdata      : out std_logic_vector(31 downto 0);                    -- readdata
			uav_writedata     : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			uav_lock          : in  std_logic                     := 'X';             -- lock
			uav_debugaccess   : in  std_logic                     := 'X';             -- debugaccess
			av_address        : out std_logic_vector(14 downto 0);                    -- address
			av_write          : out std_logic;                                        -- write
			av_readdata       : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			av_writedata      : out std_logic_vector(31 downto 0);                    -- writedata
			av_byteenable     : out std_logic_vector(3 downto 0);                     -- byteenable
			av_chipselect     : out std_logic;                                        -- chipselect
			av_clken          : out std_logic                                         -- clken
		);
	end component Nios1_onchip_memory_s1_translator;

	component Nios1_jtag_uart_avalon_jtag_slave_translator is
		port (
			clk               : in  std_logic                     := 'X';             -- clk
			reset             : in  std_logic                     := 'X';             -- reset
			uav_address       : in  std_logic_vector(18 downto 0) := (others => 'X'); -- address
			uav_burstcount    : in  std_logic_vector(2 downto 0)  := (others => 'X'); -- burstcount
			uav_read          : in  std_logic                     := 'X';             -- read
			uav_write         : in  std_logic                     := 'X';             -- write
			uav_waitrequest   : out std_logic;                                        -- waitrequest
			uav_readdatavalid : out std_logic;                                        -- readdatavalid
			uav_byteenable    : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			uav_readdata      : out std_logic_vector(31 downto 0);                    -- readdata
			uav_writedata     : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			uav_lock          : in  std_logic                     := 'X';             -- lock
			uav_debugaccess   : in  std_logic                     := 'X';             -- debugaccess
			av_address        : out std_logic;                                        -- address
			av_write          : out std_logic;                                        -- write
			av_read           : out std_logic;                                        -- read
			av_readdata       : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			av_writedata      : out std_logic_vector(31 downto 0);                    -- writedata
			av_waitrequest    : in  std_logic                     := 'X';             -- waitrequest
			av_chipselect     : out std_logic                                         -- chipselect
		);
	end component Nios1_jtag_uart_avalon_jtag_slave_translator;

	component Nios1_sysid_qsys_control_slave_translator is
		port (
			clk               : in  std_logic                     := 'X';             -- clk
			reset             : in  std_logic                     := 'X';             -- reset
			uav_address       : in  std_logic_vector(18 downto 0) := (others => 'X'); -- address
			uav_burstcount    : in  std_logic_vector(2 downto 0)  := (others => 'X'); -- burstcount
			uav_read          : in  std_logic                     := 'X';             -- read
			uav_write         : in  std_logic                     := 'X';             -- write
			uav_waitrequest   : out std_logic;                                        -- waitrequest
			uav_readdatavalid : out std_logic;                                        -- readdatavalid
			uav_byteenable    : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			uav_readdata      : out std_logic_vector(31 downto 0);                    -- readdata
			uav_writedata     : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			uav_lock          : in  std_logic                     := 'X';             -- lock
			uav_debugaccess   : in  std_logic                     := 'X';             -- debugaccess
			av_address        : out std_logic;                                        -- address
			av_readdata       : in  std_logic_vector(31 downto 0) := (others => 'X')  -- readdata
		);
	end component Nios1_sysid_qsys_control_slave_translator;

	component Nios1_pio_LEDG_s1_translator is
		port (
			clk               : in  std_logic                     := 'X';             -- clk
			reset             : in  std_logic                     := 'X';             -- reset
			uav_address       : in  std_logic_vector(18 downto 0) := (others => 'X'); -- address
			uav_burstcount    : in  std_logic_vector(2 downto 0)  := (others => 'X'); -- burstcount
			uav_read          : in  std_logic                     := 'X';             -- read
			uav_write         : in  std_logic                     := 'X';             -- write
			uav_waitrequest   : out std_logic;                                        -- waitrequest
			uav_readdatavalid : out std_logic;                                        -- readdatavalid
			uav_byteenable    : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			uav_readdata      : out std_logic_vector(31 downto 0);                    -- readdata
			uav_writedata     : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			uav_lock          : in  std_logic                     := 'X';             -- lock
			uav_debugaccess   : in  std_logic                     := 'X';             -- debugaccess
			av_address        : out std_logic_vector(2 downto 0);                     -- address
			av_write          : out std_logic;                                        -- write
			av_readdata       : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			av_writedata      : out std_logic_vector(31 downto 0);                    -- writedata
			av_chipselect     : out std_logic                                         -- chipselect
		);
	end component Nios1_pio_LEDG_s1_translator;

	component Nios1_pio_SW_s1_translator is
		port (
			clk               : in  std_logic                     := 'X';             -- clk
			reset             : in  std_logic                     := 'X';             -- reset
			uav_address       : in  std_logic_vector(18 downto 0) := (others => 'X'); -- address
			uav_burstcount    : in  std_logic_vector(2 downto 0)  := (others => 'X'); -- burstcount
			uav_read          : in  std_logic                     := 'X';             -- read
			uav_write         : in  std_logic                     := 'X';             -- write
			uav_waitrequest   : out std_logic;                                        -- waitrequest
			uav_readdatavalid : out std_logic;                                        -- readdatavalid
			uav_byteenable    : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			uav_readdata      : out std_logic_vector(31 downto 0);                    -- readdata
			uav_writedata     : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			uav_lock          : in  std_logic                     := 'X';             -- lock
			uav_debugaccess   : in  std_logic                     := 'X';             -- debugaccess
			av_address        : out std_logic_vector(1 downto 0);                     -- address
			av_readdata       : in  std_logic_vector(31 downto 0) := (others => 'X')  -- readdata
		);
	end component Nios1_pio_SW_s1_translator;

	component Nios1_pio_Button_s1_translator is
		port (
			clk               : in  std_logic                     := 'X';             -- clk
			reset             : in  std_logic                     := 'X';             -- reset
			uav_address       : in  std_logic_vector(18 downto 0) := (others => 'X'); -- address
			uav_burstcount    : in  std_logic_vector(2 downto 0)  := (others => 'X'); -- burstcount
			uav_read          : in  std_logic                     := 'X';             -- read
			uav_write         : in  std_logic                     := 'X';             -- write
			uav_waitrequest   : out std_logic;                                        -- waitrequest
			uav_readdatavalid : out std_logic;                                        -- readdatavalid
			uav_byteenable    : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			uav_readdata      : out std_logic_vector(31 downto 0);                    -- readdata
			uav_writedata     : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			uav_lock          : in  std_logic                     := 'X';             -- lock
			uav_debugaccess   : in  std_logic                     := 'X';             -- debugaccess
			av_address        : out std_logic_vector(1 downto 0);                     -- address
			av_write          : out std_logic;                                        -- write
			av_readdata       : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			av_writedata      : out std_logic_vector(31 downto 0);                    -- writedata
			av_chipselect     : out std_logic                                         -- chipselect
		);
	end component Nios1_pio_Button_s1_translator;

	component Nios1_lcd_control_slave_translator is
		port (
			clk               : in  std_logic                     := 'X';             -- clk
			reset             : in  std_logic                     := 'X';             -- reset
			uav_address       : in  std_logic_vector(18 downto 0) := (others => 'X'); -- address
			uav_burstcount    : in  std_logic_vector(2 downto 0)  := (others => 'X'); -- burstcount
			uav_read          : in  std_logic                     := 'X';             -- read
			uav_write         : in  std_logic                     := 'X';             -- write
			uav_waitrequest   : out std_logic;                                        -- waitrequest
			uav_readdatavalid : out std_logic;                                        -- readdatavalid
			uav_byteenable    : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			uav_readdata      : out std_logic_vector(31 downto 0);                    -- readdata
			uav_writedata     : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			uav_lock          : in  std_logic                     := 'X';             -- lock
			uav_debugaccess   : in  std_logic                     := 'X';             -- debugaccess
			av_address        : out std_logic_vector(1 downto 0);                     -- address
			av_write          : out std_logic;                                        -- write
			av_read           : out std_logic;                                        -- read
			av_readdata       : in  std_logic_vector(7 downto 0)  := (others => 'X'); -- readdata
			av_writedata      : out std_logic_vector(7 downto 0);                     -- writedata
			av_begintransfer  : out std_logic                                         -- begintransfer
		);
	end component Nios1_lcd_control_slave_translator;

	component Nios1_uart_s1_translator is
		port (
			clk               : in  std_logic                     := 'X';             -- clk
			reset             : in  std_logic                     := 'X';             -- reset
			uav_address       : in  std_logic_vector(18 downto 0) := (others => 'X'); -- address
			uav_burstcount    : in  std_logic_vector(2 downto 0)  := (others => 'X'); -- burstcount
			uav_read          : in  std_logic                     := 'X';             -- read
			uav_write         : in  std_logic                     := 'X';             -- write
			uav_waitrequest   : out std_logic;                                        -- waitrequest
			uav_readdatavalid : out std_logic;                                        -- readdatavalid
			uav_byteenable    : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			uav_readdata      : out std_logic_vector(31 downto 0);                    -- readdata
			uav_writedata     : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			uav_lock          : in  std_logic                     := 'X';             -- lock
			uav_debugaccess   : in  std_logic                     := 'X';             -- debugaccess
			av_address        : out std_logic_vector(2 downto 0);                     -- address
			av_write          : out std_logic;                                        -- write
			av_read           : out std_logic;                                        -- read
			av_readdata       : in  std_logic_vector(15 downto 0) := (others => 'X'); -- readdata
			av_writedata      : out std_logic_vector(15 downto 0);                    -- writedata
			av_begintransfer  : out std_logic;                                        -- begintransfer
			av_chipselect     : out std_logic                                         -- chipselect
		);
	end component Nios1_uart_s1_translator;

	component Nios1_timer_0_s1_translator is
		port (
			clk               : in  std_logic                     := 'X';             -- clk
			reset             : in  std_logic                     := 'X';             -- reset
			uav_address       : in  std_logic_vector(18 downto 0) := (others => 'X'); -- address
			uav_burstcount    : in  std_logic_vector(2 downto 0)  := (others => 'X'); -- burstcount
			uav_read          : in  std_logic                     := 'X';             -- read
			uav_write         : in  std_logic                     := 'X';             -- write
			uav_waitrequest   : out std_logic;                                        -- waitrequest
			uav_readdatavalid : out std_logic;                                        -- readdatavalid
			uav_byteenable    : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			uav_readdata      : out std_logic_vector(31 downto 0);                    -- readdata
			uav_writedata     : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			uav_lock          : in  std_logic                     := 'X';             -- lock
			uav_debugaccess   : in  std_logic                     := 'X';             -- debugaccess
			av_address        : out std_logic_vector(2 downto 0);                     -- address
			av_write          : out std_logic;                                        -- write
			av_readdata       : in  std_logic_vector(15 downto 0) := (others => 'X'); -- readdata
			av_writedata      : out std_logic_vector(15 downto 0);                    -- writedata
			av_chipselect     : out std_logic                                         -- chipselect
		);
	end component Nios1_timer_0_s1_translator;

	component Nios1_pio_LEDG_s1_translator_avalon_universal_slave_0_agent is
		port (
			clk                     : in  std_logic                     := 'X';             -- clk
			reset                   : in  std_logic                     := 'X';             -- reset
			m0_address              : out std_logic_vector(18 downto 0);                    -- address
			m0_burstcount           : out std_logic_vector(2 downto 0);                     -- burstcount
			m0_byteenable           : out std_logic_vector(3 downto 0);                     -- byteenable
			m0_debugaccess          : out std_logic;                                        -- debugaccess
			m0_lock                 : out std_logic;                                        -- lock
			m0_readdata             : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			m0_readdatavalid        : in  std_logic                     := 'X';             -- readdatavalid
			m0_read                 : out std_logic;                                        -- read
			m0_waitrequest          : in  std_logic                     := 'X';             -- waitrequest
			m0_writedata            : out std_logic_vector(31 downto 0);                    -- writedata
			m0_write                : out std_logic;                                        -- write
			rp_endofpacket          : out std_logic;                                        -- endofpacket
			rp_ready                : in  std_logic                     := 'X';             -- ready
			rp_valid                : out std_logic;                                        -- valid
			rp_data                 : out std_logic_vector(75 downto 0);                    -- data
			rp_startofpacket        : out std_logic;                                        -- startofpacket
			cp_ready                : out std_logic;                                        -- ready
			cp_valid                : in  std_logic                     := 'X';             -- valid
			cp_data                 : in  std_logic_vector(75 downto 0) := (others => 'X'); -- data
			cp_startofpacket        : in  std_logic                     := 'X';             -- startofpacket
			cp_endofpacket          : in  std_logic                     := 'X';             -- endofpacket
			cp_channel              : in  std_logic_vector(13 downto 0) := (others => 'X'); -- channel
			rf_sink_ready           : out std_logic;                                        -- ready
			rf_sink_valid           : in  std_logic                     := 'X';             -- valid
			rf_sink_startofpacket   : in  std_logic                     := 'X';             -- startofpacket
			rf_sink_endofpacket     : in  std_logic                     := 'X';             -- endofpacket
			rf_sink_data            : in  std_logic_vector(76 downto 0) := (others => 'X'); -- data
			rf_source_ready         : in  std_logic                     := 'X';             -- ready
			rf_source_valid         : out std_logic;                                        -- valid
			rf_source_startofpacket : out std_logic;                                        -- startofpacket
			rf_source_endofpacket   : out std_logic;                                        -- endofpacket
			rf_source_data          : out std_logic_vector(76 downto 0);                    -- data
			rdata_fifo_sink_ready   : out std_logic;                                        -- ready
			rdata_fifo_sink_valid   : in  std_logic                     := 'X';             -- valid
			rdata_fifo_sink_data    : in  std_logic_vector(31 downto 0) := (others => 'X'); -- data
			rdata_fifo_src_ready    : in  std_logic                     := 'X';             -- ready
			rdata_fifo_src_valid    : out std_logic;                                        -- valid
			rdata_fifo_src_data     : out std_logic_vector(31 downto 0)                     -- data
		);
	end component Nios1_pio_LEDG_s1_translator_avalon_universal_slave_0_agent;

	component Nios1_pio_LEDG_s1_translator_avalon_universal_slave_0_agent_rsp_fifo is
		port (
			clk               : in  std_logic                     := 'X';             -- clk
			reset             : in  std_logic                     := 'X';             -- reset
			in_data           : in  std_logic_vector(76 downto 0) := (others => 'X'); -- data
			in_valid          : in  std_logic                     := 'X';             -- valid
			in_ready          : out std_logic;                                        -- ready
			in_startofpacket  : in  std_logic                     := 'X';             -- startofpacket
			in_endofpacket    : in  std_logic                     := 'X';             -- endofpacket
			out_data          : out std_logic_vector(76 downto 0);                    -- data
			out_valid         : out std_logic;                                        -- valid
			out_ready         : in  std_logic                     := 'X';             -- ready
			out_startofpacket : out std_logic;                                        -- startofpacket
			out_endofpacket   : out std_logic                                         -- endofpacket
		);
	end component Nios1_pio_LEDG_s1_translator_avalon_universal_slave_0_agent_rsp_fifo;

	component Nios1_pio_LEDR_s1_translator_avalon_universal_slave_0_agent is
		port (
			clk                     : in  std_logic                     := 'X';             -- clk
			reset                   : in  std_logic                     := 'X';             -- reset
			m0_address              : out std_logic_vector(18 downto 0);                    -- address
			m0_burstcount           : out std_logic_vector(2 downto 0);                     -- burstcount
			m0_byteenable           : out std_logic_vector(3 downto 0);                     -- byteenable
			m0_debugaccess          : out std_logic;                                        -- debugaccess
			m0_lock                 : out std_logic;                                        -- lock
			m0_readdata             : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			m0_readdatavalid        : in  std_logic                     := 'X';             -- readdatavalid
			m0_read                 : out std_logic;                                        -- read
			m0_waitrequest          : in  std_logic                     := 'X';             -- waitrequest
			m0_writedata            : out std_logic_vector(31 downto 0);                    -- writedata
			m0_write                : out std_logic;                                        -- write
			rp_endofpacket          : out std_logic;                                        -- endofpacket
			rp_ready                : in  std_logic                     := 'X';             -- ready
			rp_valid                : out std_logic;                                        -- valid
			rp_data                 : out std_logic_vector(75 downto 0);                    -- data
			rp_startofpacket        : out std_logic;                                        -- startofpacket
			cp_ready                : out std_logic;                                        -- ready
			cp_valid                : in  std_logic                     := 'X';             -- valid
			cp_data                 : in  std_logic_vector(75 downto 0) := (others => 'X'); -- data
			cp_startofpacket        : in  std_logic                     := 'X';             -- startofpacket
			cp_endofpacket          : in  std_logic                     := 'X';             -- endofpacket
			cp_channel              : in  std_logic_vector(13 downto 0) := (others => 'X'); -- channel
			rf_sink_ready           : out std_logic;                                        -- ready
			rf_sink_valid           : in  std_logic                     := 'X';             -- valid
			rf_sink_startofpacket   : in  std_logic                     := 'X';             -- startofpacket
			rf_sink_endofpacket     : in  std_logic                     := 'X';             -- endofpacket
			rf_sink_data            : in  std_logic_vector(76 downto 0) := (others => 'X'); -- data
			rf_source_ready         : in  std_logic                     := 'X';             -- ready
			rf_source_valid         : out std_logic;                                        -- valid
			rf_source_startofpacket : out std_logic;                                        -- startofpacket
			rf_source_endofpacket   : out std_logic;                                        -- endofpacket
			rf_source_data          : out std_logic_vector(76 downto 0);                    -- data
			rdata_fifo_sink_ready   : out std_logic;                                        -- ready
			rdata_fifo_sink_valid   : in  std_logic                     := 'X';             -- valid
			rdata_fifo_sink_data    : in  std_logic_vector(31 downto 0) := (others => 'X'); -- data
			rdata_fifo_src_ready    : in  std_logic                     := 'X';             -- ready
			rdata_fifo_src_valid    : out std_logic;                                        -- valid
			rdata_fifo_src_data     : out std_logic_vector(31 downto 0)                     -- data
		);
	end component Nios1_pio_LEDR_s1_translator_avalon_universal_slave_0_agent;

	component Nios1_sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent is
		port (
			clk                     : in  std_logic                     := 'X';             -- clk
			reset                   : in  std_logic                     := 'X';             -- reset
			m0_address              : out std_logic_vector(18 downto 0);                    -- address
			m0_burstcount           : out std_logic_vector(2 downto 0);                     -- burstcount
			m0_byteenable           : out std_logic_vector(3 downto 0);                     -- byteenable
			m0_debugaccess          : out std_logic;                                        -- debugaccess
			m0_lock                 : out std_logic;                                        -- lock
			m0_readdata             : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			m0_readdatavalid        : in  std_logic                     := 'X';             -- readdatavalid
			m0_read                 : out std_logic;                                        -- read
			m0_waitrequest          : in  std_logic                     := 'X';             -- waitrequest
			m0_writedata            : out std_logic_vector(31 downto 0);                    -- writedata
			m0_write                : out std_logic;                                        -- write
			rp_endofpacket          : out std_logic;                                        -- endofpacket
			rp_ready                : in  std_logic                     := 'X';             -- ready
			rp_valid                : out std_logic;                                        -- valid
			rp_data                 : out std_logic_vector(75 downto 0);                    -- data
			rp_startofpacket        : out std_logic;                                        -- startofpacket
			cp_ready                : out std_logic;                                        -- ready
			cp_valid                : in  std_logic                     := 'X';             -- valid
			cp_data                 : in  std_logic_vector(75 downto 0) := (others => 'X'); -- data
			cp_startofpacket        : in  std_logic                     := 'X';             -- startofpacket
			cp_endofpacket          : in  std_logic                     := 'X';             -- endofpacket
			cp_channel              : in  std_logic_vector(13 downto 0) := (others => 'X'); -- channel
			rf_sink_ready           : out std_logic;                                        -- ready
			rf_sink_valid           : in  std_logic                     := 'X';             -- valid
			rf_sink_startofpacket   : in  std_logic                     := 'X';             -- startofpacket
			rf_sink_endofpacket     : in  std_logic                     := 'X';             -- endofpacket
			rf_sink_data            : in  std_logic_vector(76 downto 0) := (others => 'X'); -- data
			rf_source_ready         : in  std_logic                     := 'X';             -- ready
			rf_source_valid         : out std_logic;                                        -- valid
			rf_source_startofpacket : out std_logic;                                        -- startofpacket
			rf_source_endofpacket   : out std_logic;                                        -- endofpacket
			rf_source_data          : out std_logic_vector(76 downto 0);                    -- data
			rdata_fifo_sink_ready   : out std_logic;                                        -- ready
			rdata_fifo_sink_valid   : in  std_logic                     := 'X';             -- valid
			rdata_fifo_sink_data    : in  std_logic_vector(31 downto 0) := (others => 'X'); -- data
			rdata_fifo_src_ready    : in  std_logic                     := 'X';             -- ready
			rdata_fifo_src_valid    : out std_logic;                                        -- valid
			rdata_fifo_src_data     : out std_logic_vector(31 downto 0)                     -- data
		);
	end component Nios1_sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent;

	component Nios1_pio_DataRead_s1_translator_avalon_universal_slave_0_agent is
		port (
			clk                     : in  std_logic                     := 'X';             -- clk
			reset                   : in  std_logic                     := 'X';             -- reset
			m0_address              : out std_logic_vector(18 downto 0);                    -- address
			m0_burstcount           : out std_logic_vector(2 downto 0);                     -- burstcount
			m0_byteenable           : out std_logic_vector(3 downto 0);                     -- byteenable
			m0_debugaccess          : out std_logic;                                        -- debugaccess
			m0_lock                 : out std_logic;                                        -- lock
			m0_readdata             : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			m0_readdatavalid        : in  std_logic                     := 'X';             -- readdatavalid
			m0_read                 : out std_logic;                                        -- read
			m0_waitrequest          : in  std_logic                     := 'X';             -- waitrequest
			m0_writedata            : out std_logic_vector(31 downto 0);                    -- writedata
			m0_write                : out std_logic;                                        -- write
			rp_endofpacket          : out std_logic;                                        -- endofpacket
			rp_ready                : in  std_logic                     := 'X';             -- ready
			rp_valid                : out std_logic;                                        -- valid
			rp_data                 : out std_logic_vector(75 downto 0);                    -- data
			rp_startofpacket        : out std_logic;                                        -- startofpacket
			cp_ready                : out std_logic;                                        -- ready
			cp_valid                : in  std_logic                     := 'X';             -- valid
			cp_data                 : in  std_logic_vector(75 downto 0) := (others => 'X'); -- data
			cp_startofpacket        : in  std_logic                     := 'X';             -- startofpacket
			cp_endofpacket          : in  std_logic                     := 'X';             -- endofpacket
			cp_channel              : in  std_logic_vector(13 downto 0) := (others => 'X'); -- channel
			rf_sink_ready           : out std_logic;                                        -- ready
			rf_sink_valid           : in  std_logic                     := 'X';             -- valid
			rf_sink_startofpacket   : in  std_logic                     := 'X';             -- startofpacket
			rf_sink_endofpacket     : in  std_logic                     := 'X';             -- endofpacket
			rf_sink_data            : in  std_logic_vector(76 downto 0) := (others => 'X'); -- data
			rf_source_ready         : in  std_logic                     := 'X';             -- ready
			rf_source_valid         : out std_logic;                                        -- valid
			rf_source_startofpacket : out std_logic;                                        -- startofpacket
			rf_source_endofpacket   : out std_logic;                                        -- endofpacket
			rf_source_data          : out std_logic_vector(76 downto 0);                    -- data
			rdata_fifo_sink_ready   : out std_logic;                                        -- ready
			rdata_fifo_sink_valid   : in  std_logic                     := 'X';             -- valid
			rdata_fifo_sink_data    : in  std_logic_vector(31 downto 0) := (others => 'X'); -- data
			rdata_fifo_src_ready    : in  std_logic                     := 'X';             -- ready
			rdata_fifo_src_valid    : out std_logic;                                        -- valid
			rdata_fifo_src_data     : out std_logic_vector(31 downto 0)                     -- data
		);
	end component Nios1_pio_DataRead_s1_translator_avalon_universal_slave_0_agent;

	component Nios1_nios2_qsys_data_master_translator_avalon_universal_master_0_agent is
		port (
			clk              : in  std_logic                     := 'X';             -- clk
			reset            : in  std_logic                     := 'X';             -- reset
			av_address       : in  std_logic_vector(18 downto 0) := (others => 'X'); -- address
			av_write         : in  std_logic                     := 'X';             -- write
			av_read          : in  std_logic                     := 'X';             -- read
			av_writedata     : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			av_readdata      : out std_logic_vector(31 downto 0);                    -- readdata
			av_waitrequest   : out std_logic;                                        -- waitrequest
			av_readdatavalid : out std_logic;                                        -- readdatavalid
			av_byteenable    : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			av_burstcount    : in  std_logic_vector(2 downto 0)  := (others => 'X'); -- burstcount
			av_debugaccess   : in  std_logic                     := 'X';             -- debugaccess
			av_lock          : in  std_logic                     := 'X';             -- lock
			cp_valid         : out std_logic;                                        -- valid
			cp_data          : out std_logic_vector(75 downto 0);                    -- data
			cp_startofpacket : out std_logic;                                        -- startofpacket
			cp_endofpacket   : out std_logic;                                        -- endofpacket
			cp_ready         : in  std_logic                     := 'X';             -- ready
			rp_valid         : in  std_logic                     := 'X';             -- valid
			rp_data          : in  std_logic_vector(75 downto 0) := (others => 'X'); -- data
			rp_channel       : in  std_logic_vector(13 downto 0) := (others => 'X'); -- channel
			rp_startofpacket : in  std_logic                     := 'X';             -- startofpacket
			rp_endofpacket   : in  std_logic                     := 'X';             -- endofpacket
			rp_ready         : out std_logic                                         -- ready
		);
	end component Nios1_nios2_qsys_data_master_translator_avalon_universal_master_0_agent;

	component Nios1_lcd_control_slave_translator_avalon_universal_slave_0_agent is
		port (
			clk                     : in  std_logic                     := 'X';             -- clk
			reset                   : in  std_logic                     := 'X';             -- reset
			m0_address              : out std_logic_vector(18 downto 0);                    -- address
			m0_burstcount           : out std_logic_vector(2 downto 0);                     -- burstcount
			m0_byteenable           : out std_logic_vector(3 downto 0);                     -- byteenable
			m0_debugaccess          : out std_logic;                                        -- debugaccess
			m0_lock                 : out std_logic;                                        -- lock
			m0_readdata             : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			m0_readdatavalid        : in  std_logic                     := 'X';             -- readdatavalid
			m0_read                 : out std_logic;                                        -- read
			m0_waitrequest          : in  std_logic                     := 'X';             -- waitrequest
			m0_writedata            : out std_logic_vector(31 downto 0);                    -- writedata
			m0_write                : out std_logic;                                        -- write
			rp_endofpacket          : out std_logic;                                        -- endofpacket
			rp_ready                : in  std_logic                     := 'X';             -- ready
			rp_valid                : out std_logic;                                        -- valid
			rp_data                 : out std_logic_vector(75 downto 0);                    -- data
			rp_startofpacket        : out std_logic;                                        -- startofpacket
			cp_ready                : out std_logic;                                        -- ready
			cp_valid                : in  std_logic                     := 'X';             -- valid
			cp_data                 : in  std_logic_vector(75 downto 0) := (others => 'X'); -- data
			cp_startofpacket        : in  std_logic                     := 'X';             -- startofpacket
			cp_endofpacket          : in  std_logic                     := 'X';             -- endofpacket
			cp_channel              : in  std_logic_vector(13 downto 0) := (others => 'X'); -- channel
			rf_sink_ready           : out std_logic;                                        -- ready
			rf_sink_valid           : in  std_logic                     := 'X';             -- valid
			rf_sink_startofpacket   : in  std_logic                     := 'X';             -- startofpacket
			rf_sink_endofpacket     : in  std_logic                     := 'X';             -- endofpacket
			rf_sink_data            : in  std_logic_vector(76 downto 0) := (others => 'X'); -- data
			rf_source_ready         : in  std_logic                     := 'X';             -- ready
			rf_source_valid         : out std_logic;                                        -- valid
			rf_source_startofpacket : out std_logic;                                        -- startofpacket
			rf_source_endofpacket   : out std_logic;                                        -- endofpacket
			rf_source_data          : out std_logic_vector(76 downto 0);                    -- data
			rdata_fifo_sink_ready   : out std_logic;                                        -- ready
			rdata_fifo_sink_valid   : in  std_logic                     := 'X';             -- valid
			rdata_fifo_sink_data    : in  std_logic_vector(31 downto 0) := (others => 'X'); -- data
			rdata_fifo_src_ready    : in  std_logic                     := 'X';             -- ready
			rdata_fifo_src_valid    : out std_logic;                                        -- valid
			rdata_fifo_src_data     : out std_logic_vector(31 downto 0)                     -- data
		);
	end component Nios1_lcd_control_slave_translator_avalon_universal_slave_0_agent;

	component Nios1_nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent is
		port (
			clk                     : in  std_logic                     := 'X';             -- clk
			reset                   : in  std_logic                     := 'X';             -- reset
			m0_address              : out std_logic_vector(18 downto 0);                    -- address
			m0_burstcount           : out std_logic_vector(2 downto 0);                     -- burstcount
			m0_byteenable           : out std_logic_vector(3 downto 0);                     -- byteenable
			m0_debugaccess          : out std_logic;                                        -- debugaccess
			m0_lock                 : out std_logic;                                        -- lock
			m0_readdata             : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			m0_readdatavalid        : in  std_logic                     := 'X';             -- readdatavalid
			m0_read                 : out std_logic;                                        -- read
			m0_waitrequest          : in  std_logic                     := 'X';             -- waitrequest
			m0_writedata            : out std_logic_vector(31 downto 0);                    -- writedata
			m0_write                : out std_logic;                                        -- write
			rp_endofpacket          : out std_logic;                                        -- endofpacket
			rp_ready                : in  std_logic                     := 'X';             -- ready
			rp_valid                : out std_logic;                                        -- valid
			rp_data                 : out std_logic_vector(75 downto 0);                    -- data
			rp_startofpacket        : out std_logic;                                        -- startofpacket
			cp_ready                : out std_logic;                                        -- ready
			cp_valid                : in  std_logic                     := 'X';             -- valid
			cp_data                 : in  std_logic_vector(75 downto 0) := (others => 'X'); -- data
			cp_startofpacket        : in  std_logic                     := 'X';             -- startofpacket
			cp_endofpacket          : in  std_logic                     := 'X';             -- endofpacket
			cp_channel              : in  std_logic_vector(13 downto 0) := (others => 'X'); -- channel
			rf_sink_ready           : out std_logic;                                        -- ready
			rf_sink_valid           : in  std_logic                     := 'X';             -- valid
			rf_sink_startofpacket   : in  std_logic                     := 'X';             -- startofpacket
			rf_sink_endofpacket     : in  std_logic                     := 'X';             -- endofpacket
			rf_sink_data            : in  std_logic_vector(76 downto 0) := (others => 'X'); -- data
			rf_source_ready         : in  std_logic                     := 'X';             -- ready
			rf_source_valid         : out std_logic;                                        -- valid
			rf_source_startofpacket : out std_logic;                                        -- startofpacket
			rf_source_endofpacket   : out std_logic;                                        -- endofpacket
			rf_source_data          : out std_logic_vector(76 downto 0);                    -- data
			rdata_fifo_sink_ready   : out std_logic;                                        -- ready
			rdata_fifo_sink_valid   : in  std_logic                     := 'X';             -- valid
			rdata_fifo_sink_data    : in  std_logic_vector(31 downto 0) := (others => 'X'); -- data
			rdata_fifo_src_ready    : in  std_logic                     := 'X';             -- ready
			rdata_fifo_src_valid    : out std_logic;                                        -- valid
			rdata_fifo_src_data     : out std_logic_vector(31 downto 0)                     -- data
		);
	end component Nios1_nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent;

	component Nios1_nios2_qsys_instruction_master_translator_avalon_universal_master_0_agent is
		port (
			clk              : in  std_logic                     := 'X';             -- clk
			reset            : in  std_logic                     := 'X';             -- reset
			av_address       : in  std_logic_vector(18 downto 0) := (others => 'X'); -- address
			av_write         : in  std_logic                     := 'X';             -- write
			av_read          : in  std_logic                     := 'X';             -- read
			av_writedata     : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			av_readdata      : out std_logic_vector(31 downto 0);                    -- readdata
			av_waitrequest   : out std_logic;                                        -- waitrequest
			av_readdatavalid : out std_logic;                                        -- readdatavalid
			av_byteenable    : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			av_burstcount    : in  std_logic_vector(2 downto 0)  := (others => 'X'); -- burstcount
			av_debugaccess   : in  std_logic                     := 'X';             -- debugaccess
			av_lock          : in  std_logic                     := 'X';             -- lock
			cp_valid         : out std_logic;                                        -- valid
			cp_data          : out std_logic_vector(75 downto 0);                    -- data
			cp_startofpacket : out std_logic;                                        -- startofpacket
			cp_endofpacket   : out std_logic;                                        -- endofpacket
			cp_ready         : in  std_logic                     := 'X';             -- ready
			rp_valid         : in  std_logic                     := 'X';             -- valid
			rp_data          : in  std_logic_vector(75 downto 0) := (others => 'X'); -- data
			rp_channel       : in  std_logic_vector(13 downto 0) := (others => 'X'); -- channel
			rp_startofpacket : in  std_logic                     := 'X';             -- startofpacket
			rp_endofpacket   : in  std_logic                     := 'X';             -- endofpacket
			rp_ready         : out std_logic                                         -- ready
		);
	end component Nios1_nios2_qsys_instruction_master_translator_avalon_universal_master_0_agent;

	component Nios1_pio_SW_s1_translator_avalon_universal_slave_0_agent is
		port (
			clk                     : in  std_logic                     := 'X';             -- clk
			reset                   : in  std_logic                     := 'X';             -- reset
			m0_address              : out std_logic_vector(18 downto 0);                    -- address
			m0_burstcount           : out std_logic_vector(2 downto 0);                     -- burstcount
			m0_byteenable           : out std_logic_vector(3 downto 0);                     -- byteenable
			m0_debugaccess          : out std_logic;                                        -- debugaccess
			m0_lock                 : out std_logic;                                        -- lock
			m0_readdata             : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			m0_readdatavalid        : in  std_logic                     := 'X';             -- readdatavalid
			m0_read                 : out std_logic;                                        -- read
			m0_waitrequest          : in  std_logic                     := 'X';             -- waitrequest
			m0_writedata            : out std_logic_vector(31 downto 0);                    -- writedata
			m0_write                : out std_logic;                                        -- write
			rp_endofpacket          : out std_logic;                                        -- endofpacket
			rp_ready                : in  std_logic                     := 'X';             -- ready
			rp_valid                : out std_logic;                                        -- valid
			rp_data                 : out std_logic_vector(75 downto 0);                    -- data
			rp_startofpacket        : out std_logic;                                        -- startofpacket
			cp_ready                : out std_logic;                                        -- ready
			cp_valid                : in  std_logic                     := 'X';             -- valid
			cp_data                 : in  std_logic_vector(75 downto 0) := (others => 'X'); -- data
			cp_startofpacket        : in  std_logic                     := 'X';             -- startofpacket
			cp_endofpacket          : in  std_logic                     := 'X';             -- endofpacket
			cp_channel              : in  std_logic_vector(13 downto 0) := (others => 'X'); -- channel
			rf_sink_ready           : out std_logic;                                        -- ready
			rf_sink_valid           : in  std_logic                     := 'X';             -- valid
			rf_sink_startofpacket   : in  std_logic                     := 'X';             -- startofpacket
			rf_sink_endofpacket     : in  std_logic                     := 'X';             -- endofpacket
			rf_sink_data            : in  std_logic_vector(76 downto 0) := (others => 'X'); -- data
			rf_source_ready         : in  std_logic                     := 'X';             -- ready
			rf_source_valid         : out std_logic;                                        -- valid
			rf_source_startofpacket : out std_logic;                                        -- startofpacket
			rf_source_endofpacket   : out std_logic;                                        -- endofpacket
			rf_source_data          : out std_logic_vector(76 downto 0);                    -- data
			rdata_fifo_sink_ready   : out std_logic;                                        -- ready
			rdata_fifo_sink_valid   : in  std_logic                     := 'X';             -- valid
			rdata_fifo_sink_data    : in  std_logic_vector(31 downto 0) := (others => 'X'); -- data
			rdata_fifo_src_ready    : in  std_logic                     := 'X';             -- ready
			rdata_fifo_src_valid    : out std_logic;                                        -- valid
			rdata_fifo_src_data     : out std_logic_vector(31 downto 0)                     -- data
		);
	end component Nios1_pio_SW_s1_translator_avalon_universal_slave_0_agent;

	component Nios1_jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent is
		port (
			clk                     : in  std_logic                     := 'X';             -- clk
			reset                   : in  std_logic                     := 'X';             -- reset
			m0_address              : out std_logic_vector(18 downto 0);                    -- address
			m0_burstcount           : out std_logic_vector(2 downto 0);                     -- burstcount
			m0_byteenable           : out std_logic_vector(3 downto 0);                     -- byteenable
			m0_debugaccess          : out std_logic;                                        -- debugaccess
			m0_lock                 : out std_logic;                                        -- lock
			m0_readdata             : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			m0_readdatavalid        : in  std_logic                     := 'X';             -- readdatavalid
			m0_read                 : out std_logic;                                        -- read
			m0_waitrequest          : in  std_logic                     := 'X';             -- waitrequest
			m0_writedata            : out std_logic_vector(31 downto 0);                    -- writedata
			m0_write                : out std_logic;                                        -- write
			rp_endofpacket          : out std_logic;                                        -- endofpacket
			rp_ready                : in  std_logic                     := 'X';             -- ready
			rp_valid                : out std_logic;                                        -- valid
			rp_data                 : out std_logic_vector(75 downto 0);                    -- data
			rp_startofpacket        : out std_logic;                                        -- startofpacket
			cp_ready                : out std_logic;                                        -- ready
			cp_valid                : in  std_logic                     := 'X';             -- valid
			cp_data                 : in  std_logic_vector(75 downto 0) := (others => 'X'); -- data
			cp_startofpacket        : in  std_logic                     := 'X';             -- startofpacket
			cp_endofpacket          : in  std_logic                     := 'X';             -- endofpacket
			cp_channel              : in  std_logic_vector(13 downto 0) := (others => 'X'); -- channel
			rf_sink_ready           : out std_logic;                                        -- ready
			rf_sink_valid           : in  std_logic                     := 'X';             -- valid
			rf_sink_startofpacket   : in  std_logic                     := 'X';             -- startofpacket
			rf_sink_endofpacket     : in  std_logic                     := 'X';             -- endofpacket
			rf_sink_data            : in  std_logic_vector(76 downto 0) := (others => 'X'); -- data
			rf_source_ready         : in  std_logic                     := 'X';             -- ready
			rf_source_valid         : out std_logic;                                        -- valid
			rf_source_startofpacket : out std_logic;                                        -- startofpacket
			rf_source_endofpacket   : out std_logic;                                        -- endofpacket
			rf_source_data          : out std_logic_vector(76 downto 0);                    -- data
			rdata_fifo_sink_ready   : out std_logic;                                        -- ready
			rdata_fifo_sink_valid   : in  std_logic                     := 'X';             -- valid
			rdata_fifo_sink_data    : in  std_logic_vector(31 downto 0) := (others => 'X'); -- data
			rdata_fifo_src_ready    : in  std_logic                     := 'X';             -- ready
			rdata_fifo_src_valid    : out std_logic;                                        -- valid
			rdata_fifo_src_data     : out std_logic_vector(31 downto 0)                     -- data
		);
	end component Nios1_jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent;

	component Nios1_pio_Button_s1_translator_avalon_universal_slave_0_agent is
		port (
			clk                     : in  std_logic                     := 'X';             -- clk
			reset                   : in  std_logic                     := 'X';             -- reset
			m0_address              : out std_logic_vector(18 downto 0);                    -- address
			m0_burstcount           : out std_logic_vector(2 downto 0);                     -- burstcount
			m0_byteenable           : out std_logic_vector(3 downto 0);                     -- byteenable
			m0_debugaccess          : out std_logic;                                        -- debugaccess
			m0_lock                 : out std_logic;                                        -- lock
			m0_readdata             : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			m0_readdatavalid        : in  std_logic                     := 'X';             -- readdatavalid
			m0_read                 : out std_logic;                                        -- read
			m0_waitrequest          : in  std_logic                     := 'X';             -- waitrequest
			m0_writedata            : out std_logic_vector(31 downto 0);                    -- writedata
			m0_write                : out std_logic;                                        -- write
			rp_endofpacket          : out std_logic;                                        -- endofpacket
			rp_ready                : in  std_logic                     := 'X';             -- ready
			rp_valid                : out std_logic;                                        -- valid
			rp_data                 : out std_logic_vector(75 downto 0);                    -- data
			rp_startofpacket        : out std_logic;                                        -- startofpacket
			cp_ready                : out std_logic;                                        -- ready
			cp_valid                : in  std_logic                     := 'X';             -- valid
			cp_data                 : in  std_logic_vector(75 downto 0) := (others => 'X'); -- data
			cp_startofpacket        : in  std_logic                     := 'X';             -- startofpacket
			cp_endofpacket          : in  std_logic                     := 'X';             -- endofpacket
			cp_channel              : in  std_logic_vector(13 downto 0) := (others => 'X'); -- channel
			rf_sink_ready           : out std_logic;                                        -- ready
			rf_sink_valid           : in  std_logic                     := 'X';             -- valid
			rf_sink_startofpacket   : in  std_logic                     := 'X';             -- startofpacket
			rf_sink_endofpacket     : in  std_logic                     := 'X';             -- endofpacket
			rf_sink_data            : in  std_logic_vector(76 downto 0) := (others => 'X'); -- data
			rf_source_ready         : in  std_logic                     := 'X';             -- ready
			rf_source_valid         : out std_logic;                                        -- valid
			rf_source_startofpacket : out std_logic;                                        -- startofpacket
			rf_source_endofpacket   : out std_logic;                                        -- endofpacket
			rf_source_data          : out std_logic_vector(76 downto 0);                    -- data
			rdata_fifo_sink_ready   : out std_logic;                                        -- ready
			rdata_fifo_sink_valid   : in  std_logic                     := 'X';             -- valid
			rdata_fifo_sink_data    : in  std_logic_vector(31 downto 0) := (others => 'X'); -- data
			rdata_fifo_src_ready    : in  std_logic                     := 'X';             -- ready
			rdata_fifo_src_valid    : out std_logic;                                        -- valid
			rdata_fifo_src_data     : out std_logic_vector(31 downto 0)                     -- data
		);
	end component Nios1_pio_Button_s1_translator_avalon_universal_slave_0_agent;

	component Nios1_pio_Data_s1_translator_avalon_universal_slave_0_agent is
		port (
			clk                     : in  std_logic                     := 'X';             -- clk
			reset                   : in  std_logic                     := 'X';             -- reset
			m0_address              : out std_logic_vector(18 downto 0);                    -- address
			m0_burstcount           : out std_logic_vector(2 downto 0);                     -- burstcount
			m0_byteenable           : out std_logic_vector(3 downto 0);                     -- byteenable
			m0_debugaccess          : out std_logic;                                        -- debugaccess
			m0_lock                 : out std_logic;                                        -- lock
			m0_readdata             : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			m0_readdatavalid        : in  std_logic                     := 'X';             -- readdatavalid
			m0_read                 : out std_logic;                                        -- read
			m0_waitrequest          : in  std_logic                     := 'X';             -- waitrequest
			m0_writedata            : out std_logic_vector(31 downto 0);                    -- writedata
			m0_write                : out std_logic;                                        -- write
			rp_endofpacket          : out std_logic;                                        -- endofpacket
			rp_ready                : in  std_logic                     := 'X';             -- ready
			rp_valid                : out std_logic;                                        -- valid
			rp_data                 : out std_logic_vector(75 downto 0);                    -- data
			rp_startofpacket        : out std_logic;                                        -- startofpacket
			cp_ready                : out std_logic;                                        -- ready
			cp_valid                : in  std_logic                     := 'X';             -- valid
			cp_data                 : in  std_logic_vector(75 downto 0) := (others => 'X'); -- data
			cp_startofpacket        : in  std_logic                     := 'X';             -- startofpacket
			cp_endofpacket          : in  std_logic                     := 'X';             -- endofpacket
			cp_channel              : in  std_logic_vector(13 downto 0) := (others => 'X'); -- channel
			rf_sink_ready           : out std_logic;                                        -- ready
			rf_sink_valid           : in  std_logic                     := 'X';             -- valid
			rf_sink_startofpacket   : in  std_logic                     := 'X';             -- startofpacket
			rf_sink_endofpacket     : in  std_logic                     := 'X';             -- endofpacket
			rf_sink_data            : in  std_logic_vector(76 downto 0) := (others => 'X'); -- data
			rf_source_ready         : in  std_logic                     := 'X';             -- ready
			rf_source_valid         : out std_logic;                                        -- valid
			rf_source_startofpacket : out std_logic;                                        -- startofpacket
			rf_source_endofpacket   : out std_logic;                                        -- endofpacket
			rf_source_data          : out std_logic_vector(76 downto 0);                    -- data
			rdata_fifo_sink_ready   : out std_logic;                                        -- ready
			rdata_fifo_sink_valid   : in  std_logic                     := 'X';             -- valid
			rdata_fifo_sink_data    : in  std_logic_vector(31 downto 0) := (others => 'X'); -- data
			rdata_fifo_src_ready    : in  std_logic                     := 'X';             -- ready
			rdata_fifo_src_valid    : out std_logic;                                        -- valid
			rdata_fifo_src_data     : out std_logic_vector(31 downto 0)                     -- data
		);
	end component Nios1_pio_Data_s1_translator_avalon_universal_slave_0_agent;

	component Nios1_uart_s1_translator_avalon_universal_slave_0_agent is
		port (
			clk                     : in  std_logic                     := 'X';             -- clk
			reset                   : in  std_logic                     := 'X';             -- reset
			m0_address              : out std_logic_vector(18 downto 0);                    -- address
			m0_burstcount           : out std_logic_vector(2 downto 0);                     -- burstcount
			m0_byteenable           : out std_logic_vector(3 downto 0);                     -- byteenable
			m0_debugaccess          : out std_logic;                                        -- debugaccess
			m0_lock                 : out std_logic;                                        -- lock
			m0_readdata             : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			m0_readdatavalid        : in  std_logic                     := 'X';             -- readdatavalid
			m0_read                 : out std_logic;                                        -- read
			m0_waitrequest          : in  std_logic                     := 'X';             -- waitrequest
			m0_writedata            : out std_logic_vector(31 downto 0);                    -- writedata
			m0_write                : out std_logic;                                        -- write
			rp_endofpacket          : out std_logic;                                        -- endofpacket
			rp_ready                : in  std_logic                     := 'X';             -- ready
			rp_valid                : out std_logic;                                        -- valid
			rp_data                 : out std_logic_vector(75 downto 0);                    -- data
			rp_startofpacket        : out std_logic;                                        -- startofpacket
			cp_ready                : out std_logic;                                        -- ready
			cp_valid                : in  std_logic                     := 'X';             -- valid
			cp_data                 : in  std_logic_vector(75 downto 0) := (others => 'X'); -- data
			cp_startofpacket        : in  std_logic                     := 'X';             -- startofpacket
			cp_endofpacket          : in  std_logic                     := 'X';             -- endofpacket
			cp_channel              : in  std_logic_vector(13 downto 0) := (others => 'X'); -- channel
			rf_sink_ready           : out std_logic;                                        -- ready
			rf_sink_valid           : in  std_logic                     := 'X';             -- valid
			rf_sink_startofpacket   : in  std_logic                     := 'X';             -- startofpacket
			rf_sink_endofpacket     : in  std_logic                     := 'X';             -- endofpacket
			rf_sink_data            : in  std_logic_vector(76 downto 0) := (others => 'X'); -- data
			rf_source_ready         : in  std_logic                     := 'X';             -- ready
			rf_source_valid         : out std_logic;                                        -- valid
			rf_source_startofpacket : out std_logic;                                        -- startofpacket
			rf_source_endofpacket   : out std_logic;                                        -- endofpacket
			rf_source_data          : out std_logic_vector(76 downto 0);                    -- data
			rdata_fifo_sink_ready   : out std_logic;                                        -- ready
			rdata_fifo_sink_valid   : in  std_logic                     := 'X';             -- valid
			rdata_fifo_sink_data    : in  std_logic_vector(31 downto 0) := (others => 'X'); -- data
			rdata_fifo_src_ready    : in  std_logic                     := 'X';             -- ready
			rdata_fifo_src_valid    : out std_logic;                                        -- valid
			rdata_fifo_src_data     : out std_logic_vector(31 downto 0)                     -- data
		);
	end component Nios1_uart_s1_translator_avalon_universal_slave_0_agent;

	component Nios1_onchip_memory_s1_translator_avalon_universal_slave_0_agent is
		port (
			clk                     : in  std_logic                     := 'X';             -- clk
			reset                   : in  std_logic                     := 'X';             -- reset
			m0_address              : out std_logic_vector(18 downto 0);                    -- address
			m0_burstcount           : out std_logic_vector(2 downto 0);                     -- burstcount
			m0_byteenable           : out std_logic_vector(3 downto 0);                     -- byteenable
			m0_debugaccess          : out std_logic;                                        -- debugaccess
			m0_lock                 : out std_logic;                                        -- lock
			m0_readdata             : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			m0_readdatavalid        : in  std_logic                     := 'X';             -- readdatavalid
			m0_read                 : out std_logic;                                        -- read
			m0_waitrequest          : in  std_logic                     := 'X';             -- waitrequest
			m0_writedata            : out std_logic_vector(31 downto 0);                    -- writedata
			m0_write                : out std_logic;                                        -- write
			rp_endofpacket          : out std_logic;                                        -- endofpacket
			rp_ready                : in  std_logic                     := 'X';             -- ready
			rp_valid                : out std_logic;                                        -- valid
			rp_data                 : out std_logic_vector(75 downto 0);                    -- data
			rp_startofpacket        : out std_logic;                                        -- startofpacket
			cp_ready                : out std_logic;                                        -- ready
			cp_valid                : in  std_logic                     := 'X';             -- valid
			cp_data                 : in  std_logic_vector(75 downto 0) := (others => 'X'); -- data
			cp_startofpacket        : in  std_logic                     := 'X';             -- startofpacket
			cp_endofpacket          : in  std_logic                     := 'X';             -- endofpacket
			cp_channel              : in  std_logic_vector(13 downto 0) := (others => 'X'); -- channel
			rf_sink_ready           : out std_logic;                                        -- ready
			rf_sink_valid           : in  std_logic                     := 'X';             -- valid
			rf_sink_startofpacket   : in  std_logic                     := 'X';             -- startofpacket
			rf_sink_endofpacket     : in  std_logic                     := 'X';             -- endofpacket
			rf_sink_data            : in  std_logic_vector(76 downto 0) := (others => 'X'); -- data
			rf_source_ready         : in  std_logic                     := 'X';             -- ready
			rf_source_valid         : out std_logic;                                        -- valid
			rf_source_startofpacket : out std_logic;                                        -- startofpacket
			rf_source_endofpacket   : out std_logic;                                        -- endofpacket
			rf_source_data          : out std_logic_vector(76 downto 0);                    -- data
			rdata_fifo_sink_ready   : out std_logic;                                        -- ready
			rdata_fifo_sink_valid   : in  std_logic                     := 'X';             -- valid
			rdata_fifo_sink_data    : in  std_logic_vector(31 downto 0) := (others => 'X'); -- data
			rdata_fifo_src_ready    : in  std_logic                     := 'X';             -- ready
			rdata_fifo_src_valid    : out std_logic;                                        -- valid
			rdata_fifo_src_data     : out std_logic_vector(31 downto 0)                     -- data
		);
	end component Nios1_onchip_memory_s1_translator_avalon_universal_slave_0_agent;

	component Nios1_timer_0_s1_translator_avalon_universal_slave_0_agent is
		port (
			clk                     : in  std_logic                     := 'X';             -- clk
			reset                   : in  std_logic                     := 'X';             -- reset
			m0_address              : out std_logic_vector(18 downto 0);                    -- address
			m0_burstcount           : out std_logic_vector(2 downto 0);                     -- burstcount
			m0_byteenable           : out std_logic_vector(3 downto 0);                     -- byteenable
			m0_debugaccess          : out std_logic;                                        -- debugaccess
			m0_lock                 : out std_logic;                                        -- lock
			m0_readdata             : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			m0_readdatavalid        : in  std_logic                     := 'X';             -- readdatavalid
			m0_read                 : out std_logic;                                        -- read
			m0_waitrequest          : in  std_logic                     := 'X';             -- waitrequest
			m0_writedata            : out std_logic_vector(31 downto 0);                    -- writedata
			m0_write                : out std_logic;                                        -- write
			rp_endofpacket          : out std_logic;                                        -- endofpacket
			rp_ready                : in  std_logic                     := 'X';             -- ready
			rp_valid                : out std_logic;                                        -- valid
			rp_data                 : out std_logic_vector(75 downto 0);                    -- data
			rp_startofpacket        : out std_logic;                                        -- startofpacket
			cp_ready                : out std_logic;                                        -- ready
			cp_valid                : in  std_logic                     := 'X';             -- valid
			cp_data                 : in  std_logic_vector(75 downto 0) := (others => 'X'); -- data
			cp_startofpacket        : in  std_logic                     := 'X';             -- startofpacket
			cp_endofpacket          : in  std_logic                     := 'X';             -- endofpacket
			cp_channel              : in  std_logic_vector(13 downto 0) := (others => 'X'); -- channel
			rf_sink_ready           : out std_logic;                                        -- ready
			rf_sink_valid           : in  std_logic                     := 'X';             -- valid
			rf_sink_startofpacket   : in  std_logic                     := 'X';             -- startofpacket
			rf_sink_endofpacket     : in  std_logic                     := 'X';             -- endofpacket
			rf_sink_data            : in  std_logic_vector(76 downto 0) := (others => 'X'); -- data
			rf_source_ready         : in  std_logic                     := 'X';             -- ready
			rf_source_valid         : out std_logic;                                        -- valid
			rf_source_startofpacket : out std_logic;                                        -- startofpacket
			rf_source_endofpacket   : out std_logic;                                        -- endofpacket
			rf_source_data          : out std_logic_vector(76 downto 0);                    -- data
			rdata_fifo_sink_ready   : out std_logic;                                        -- ready
			rdata_fifo_sink_valid   : in  std_logic                     := 'X';             -- valid
			rdata_fifo_sink_data    : in  std_logic_vector(31 downto 0) := (others => 'X'); -- data
			rdata_fifo_src_ready    : in  std_logic                     := 'X';             -- ready
			rdata_fifo_src_valid    : out std_logic;                                        -- valid
			rdata_fifo_src_data     : out std_logic_vector(31 downto 0)                     -- data
		);
	end component Nios1_timer_0_s1_translator_avalon_universal_slave_0_agent;

	component Nios1_pio_RdyData_s1_translator_avalon_universal_slave_0_agent is
		port (
			clk                     : in  std_logic                     := 'X';             -- clk
			reset                   : in  std_logic                     := 'X';             -- reset
			m0_address              : out std_logic_vector(18 downto 0);                    -- address
			m0_burstcount           : out std_logic_vector(2 downto 0);                     -- burstcount
			m0_byteenable           : out std_logic_vector(3 downto 0);                     -- byteenable
			m0_debugaccess          : out std_logic;                                        -- debugaccess
			m0_lock                 : out std_logic;                                        -- lock
			m0_readdata             : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			m0_readdatavalid        : in  std_logic                     := 'X';             -- readdatavalid
			m0_read                 : out std_logic;                                        -- read
			m0_waitrequest          : in  std_logic                     := 'X';             -- waitrequest
			m0_writedata            : out std_logic_vector(31 downto 0);                    -- writedata
			m0_write                : out std_logic;                                        -- write
			rp_endofpacket          : out std_logic;                                        -- endofpacket
			rp_ready                : in  std_logic                     := 'X';             -- ready
			rp_valid                : out std_logic;                                        -- valid
			rp_data                 : out std_logic_vector(75 downto 0);                    -- data
			rp_startofpacket        : out std_logic;                                        -- startofpacket
			cp_ready                : out std_logic;                                        -- ready
			cp_valid                : in  std_logic                     := 'X';             -- valid
			cp_data                 : in  std_logic_vector(75 downto 0) := (others => 'X'); -- data
			cp_startofpacket        : in  std_logic                     := 'X';             -- startofpacket
			cp_endofpacket          : in  std_logic                     := 'X';             -- endofpacket
			cp_channel              : in  std_logic_vector(13 downto 0) := (others => 'X'); -- channel
			rf_sink_ready           : out std_logic;                                        -- ready
			rf_sink_valid           : in  std_logic                     := 'X';             -- valid
			rf_sink_startofpacket   : in  std_logic                     := 'X';             -- startofpacket
			rf_sink_endofpacket     : in  std_logic                     := 'X';             -- endofpacket
			rf_sink_data            : in  std_logic_vector(76 downto 0) := (others => 'X'); -- data
			rf_source_ready         : in  std_logic                     := 'X';             -- ready
			rf_source_valid         : out std_logic;                                        -- valid
			rf_source_startofpacket : out std_logic;                                        -- startofpacket
			rf_source_endofpacket   : out std_logic;                                        -- endofpacket
			rf_source_data          : out std_logic_vector(76 downto 0);                    -- data
			rdata_fifo_sink_ready   : out std_logic;                                        -- ready
			rdata_fifo_sink_valid   : in  std_logic                     := 'X';             -- valid
			rdata_fifo_sink_data    : in  std_logic_vector(31 downto 0) := (others => 'X'); -- data
			rdata_fifo_src_ready    : in  std_logic                     := 'X';             -- ready
			rdata_fifo_src_valid    : out std_logic;                                        -- valid
			rdata_fifo_src_data     : out std_logic_vector(31 downto 0)                     -- data
		);
	end component Nios1_pio_RdyData_s1_translator_avalon_universal_slave_0_agent;

	component Nios1_addr_router is
		port (
			sink_ready         : out std_logic;                                        -- ready
			sink_valid         : in  std_logic                     := 'X';             -- valid
			sink_data          : in  std_logic_vector(75 downto 0) := (others => 'X'); -- data
			sink_startofpacket : in  std_logic                     := 'X';             -- startofpacket
			sink_endofpacket   : in  std_logic                     := 'X';             -- endofpacket
			clk                : in  std_logic                     := 'X';             -- clk
			reset              : in  std_logic                     := 'X';             -- reset
			src_ready          : in  std_logic                     := 'X';             -- ready
			src_valid          : out std_logic;                                        -- valid
			src_data           : out std_logic_vector(75 downto 0);                    -- data
			src_channel        : out std_logic_vector(13 downto 0);                    -- channel
			src_startofpacket  : out std_logic;                                        -- startofpacket
			src_endofpacket    : out std_logic                                         -- endofpacket
		);
	end component Nios1_addr_router;

	component Nios1_addr_router_001 is
		port (
			sink_ready         : out std_logic;                                        -- ready
			sink_valid         : in  std_logic                     := 'X';             -- valid
			sink_data          : in  std_logic_vector(75 downto 0) := (others => 'X'); -- data
			sink_startofpacket : in  std_logic                     := 'X';             -- startofpacket
			sink_endofpacket   : in  std_logic                     := 'X';             -- endofpacket
			clk                : in  std_logic                     := 'X';             -- clk
			reset              : in  std_logic                     := 'X';             -- reset
			src_ready          : in  std_logic                     := 'X';             -- ready
			src_valid          : out std_logic;                                        -- valid
			src_data           : out std_logic_vector(75 downto 0);                    -- data
			src_channel        : out std_logic_vector(13 downto 0);                    -- channel
			src_startofpacket  : out std_logic;                                        -- startofpacket
			src_endofpacket    : out std_logic                                         -- endofpacket
		);
	end component Nios1_addr_router_001;

	component Nios1_id_router is
		port (
			sink_ready         : out std_logic;                                        -- ready
			sink_valid         : in  std_logic                     := 'X';             -- valid
			sink_data          : in  std_logic_vector(75 downto 0) := (others => 'X'); -- data
			sink_startofpacket : in  std_logic                     := 'X';             -- startofpacket
			sink_endofpacket   : in  std_logic                     := 'X';             -- endofpacket
			clk                : in  std_logic                     := 'X';             -- clk
			reset              : in  std_logic                     := 'X';             -- reset
			src_ready          : in  std_logic                     := 'X';             -- ready
			src_valid          : out std_logic;                                        -- valid
			src_data           : out std_logic_vector(75 downto 0);                    -- data
			src_channel        : out std_logic_vector(13 downto 0);                    -- channel
			src_startofpacket  : out std_logic;                                        -- startofpacket
			src_endofpacket    : out std_logic                                         -- endofpacket
		);
	end component Nios1_id_router;

	component Nios1_id_router_002 is
		port (
			sink_ready         : out std_logic;                                        -- ready
			sink_valid         : in  std_logic                     := 'X';             -- valid
			sink_data          : in  std_logic_vector(75 downto 0) := (others => 'X'); -- data
			sink_startofpacket : in  std_logic                     := 'X';             -- startofpacket
			sink_endofpacket   : in  std_logic                     := 'X';             -- endofpacket
			clk                : in  std_logic                     := 'X';             -- clk
			reset              : in  std_logic                     := 'X';             -- reset
			src_ready          : in  std_logic                     := 'X';             -- ready
			src_valid          : out std_logic;                                        -- valid
			src_data           : out std_logic_vector(75 downto 0);                    -- data
			src_channel        : out std_logic_vector(13 downto 0);                    -- channel
			src_startofpacket  : out std_logic;                                        -- startofpacket
			src_endofpacket    : out std_logic                                         -- endofpacket
		);
	end component Nios1_id_router_002;

	component Nios1_limiter is
		port (
			clk                    : in  std_logic                     := 'X';             -- clk
			reset                  : in  std_logic                     := 'X';             -- reset
			cmd_sink_ready         : out std_logic;                                        -- ready
			cmd_sink_valid         : in  std_logic                     := 'X';             -- valid
			cmd_sink_data          : in  std_logic_vector(75 downto 0) := (others => 'X'); -- data
			cmd_sink_channel       : in  std_logic_vector(13 downto 0) := (others => 'X'); -- channel
			cmd_sink_startofpacket : in  std_logic                     := 'X';             -- startofpacket
			cmd_sink_endofpacket   : in  std_logic                     := 'X';             -- endofpacket
			cmd_src_ready          : in  std_logic                     := 'X';             -- ready
			cmd_src_data           : out std_logic_vector(75 downto 0);                    -- data
			cmd_src_channel        : out std_logic_vector(13 downto 0);                    -- channel
			cmd_src_startofpacket  : out std_logic;                                        -- startofpacket
			cmd_src_endofpacket    : out std_logic;                                        -- endofpacket
			rsp_sink_ready         : out std_logic;                                        -- ready
			rsp_sink_valid         : in  std_logic                     := 'X';             -- valid
			rsp_sink_channel       : in  std_logic_vector(13 downto 0) := (others => 'X'); -- channel
			rsp_sink_data          : in  std_logic_vector(75 downto 0) := (others => 'X'); -- data
			rsp_sink_startofpacket : in  std_logic                     := 'X';             -- startofpacket
			rsp_sink_endofpacket   : in  std_logic                     := 'X';             -- endofpacket
			rsp_src_ready          : in  std_logic                     := 'X';             -- ready
			rsp_src_valid          : out std_logic;                                        -- valid
			rsp_src_data           : out std_logic_vector(75 downto 0);                    -- data
			rsp_src_channel        : out std_logic_vector(13 downto 0);                    -- channel
			rsp_src_startofpacket  : out std_logic;                                        -- startofpacket
			rsp_src_endofpacket    : out std_logic;                                        -- endofpacket
			cmd_src_valid          : out std_logic_vector(13 downto 0)                     -- data
		);
	end component Nios1_limiter;

	component Nios1_rst_controller is
		port (
			reset_in0 : in  std_logic := 'X'; -- reset
			clk       : in  std_logic := 'X'; -- clk
			reset_out : out std_logic         -- reset
		);
	end component Nios1_rst_controller;

	component Nios1_cmd_xbar_demux is
		port (
			clk                : in  std_logic                     := 'X';             -- clk
			reset              : in  std_logic                     := 'X';             -- reset
			sink_ready         : out std_logic;                                        -- ready
			sink_channel       : in  std_logic_vector(13 downto 0) := (others => 'X'); -- channel
			sink_data          : in  std_logic_vector(75 downto 0) := (others => 'X'); -- data
			sink_startofpacket : in  std_logic                     := 'X';             -- startofpacket
			sink_endofpacket   : in  std_logic                     := 'X';             -- endofpacket
			sink_valid         : in  std_logic_vector(13 downto 0) := (others => 'X'); -- data
			src0_ready         : in  std_logic                     := 'X';             -- ready
			src0_valid         : out std_logic;                                        -- valid
			src0_data          : out std_logic_vector(75 downto 0);                    -- data
			src0_channel       : out std_logic_vector(13 downto 0);                    -- channel
			src0_startofpacket : out std_logic;                                        -- startofpacket
			src0_endofpacket   : out std_logic;                                        -- endofpacket
			src1_ready         : in  std_logic                     := 'X';             -- ready
			src1_valid         : out std_logic;                                        -- valid
			src1_data          : out std_logic_vector(75 downto 0);                    -- data
			src1_channel       : out std_logic_vector(13 downto 0);                    -- channel
			src1_startofpacket : out std_logic;                                        -- startofpacket
			src1_endofpacket   : out std_logic                                         -- endofpacket
		);
	end component Nios1_cmd_xbar_demux;

	component Nios1_cmd_xbar_demux_001 is
		port (
			clk                 : in  std_logic                     := 'X';             -- clk
			reset               : in  std_logic                     := 'X';             -- reset
			sink_ready          : out std_logic;                                        -- ready
			sink_channel        : in  std_logic_vector(13 downto 0) := (others => 'X'); -- channel
			sink_data           : in  std_logic_vector(75 downto 0) := (others => 'X'); -- data
			sink_startofpacket  : in  std_logic                     := 'X';             -- startofpacket
			sink_endofpacket    : in  std_logic                     := 'X';             -- endofpacket
			sink_valid          : in  std_logic_vector(13 downto 0) := (others => 'X'); -- data
			src0_ready          : in  std_logic                     := 'X';             -- ready
			src0_valid          : out std_logic;                                        -- valid
			src0_data           : out std_logic_vector(75 downto 0);                    -- data
			src0_channel        : out std_logic_vector(13 downto 0);                    -- channel
			src0_startofpacket  : out std_logic;                                        -- startofpacket
			src0_endofpacket    : out std_logic;                                        -- endofpacket
			src1_ready          : in  std_logic                     := 'X';             -- ready
			src1_valid          : out std_logic;                                        -- valid
			src1_data           : out std_logic_vector(75 downto 0);                    -- data
			src1_channel        : out std_logic_vector(13 downto 0);                    -- channel
			src1_startofpacket  : out std_logic;                                        -- startofpacket
			src1_endofpacket    : out std_logic;                                        -- endofpacket
			src2_ready          : in  std_logic                     := 'X';             -- ready
			src2_valid          : out std_logic;                                        -- valid
			src2_data           : out std_logic_vector(75 downto 0);                    -- data
			src2_channel        : out std_logic_vector(13 downto 0);                    -- channel
			src2_startofpacket  : out std_logic;                                        -- startofpacket
			src2_endofpacket    : out std_logic;                                        -- endofpacket
			src3_ready          : in  std_logic                     := 'X';             -- ready
			src3_valid          : out std_logic;                                        -- valid
			src3_data           : out std_logic_vector(75 downto 0);                    -- data
			src3_channel        : out std_logic_vector(13 downto 0);                    -- channel
			src3_startofpacket  : out std_logic;                                        -- startofpacket
			src3_endofpacket    : out std_logic;                                        -- endofpacket
			src4_ready          : in  std_logic                     := 'X';             -- ready
			src4_valid          : out std_logic;                                        -- valid
			src4_data           : out std_logic_vector(75 downto 0);                    -- data
			src4_channel        : out std_logic_vector(13 downto 0);                    -- channel
			src4_startofpacket  : out std_logic;                                        -- startofpacket
			src4_endofpacket    : out std_logic;                                        -- endofpacket
			src5_ready          : in  std_logic                     := 'X';             -- ready
			src5_valid          : out std_logic;                                        -- valid
			src5_data           : out std_logic_vector(75 downto 0);                    -- data
			src5_channel        : out std_logic_vector(13 downto 0);                    -- channel
			src5_startofpacket  : out std_logic;                                        -- startofpacket
			src5_endofpacket    : out std_logic;                                        -- endofpacket
			src6_ready          : in  std_logic                     := 'X';             -- ready
			src6_valid          : out std_logic;                                        -- valid
			src6_data           : out std_logic_vector(75 downto 0);                    -- data
			src6_channel        : out std_logic_vector(13 downto 0);                    -- channel
			src6_startofpacket  : out std_logic;                                        -- startofpacket
			src6_endofpacket    : out std_logic;                                        -- endofpacket
			src7_ready          : in  std_logic                     := 'X';             -- ready
			src7_valid          : out std_logic;                                        -- valid
			src7_data           : out std_logic_vector(75 downto 0);                    -- data
			src7_channel        : out std_logic_vector(13 downto 0);                    -- channel
			src7_startofpacket  : out std_logic;                                        -- startofpacket
			src7_endofpacket    : out std_logic;                                        -- endofpacket
			src8_ready          : in  std_logic                     := 'X';             -- ready
			src8_valid          : out std_logic;                                        -- valid
			src8_data           : out std_logic_vector(75 downto 0);                    -- data
			src8_channel        : out std_logic_vector(13 downto 0);                    -- channel
			src8_startofpacket  : out std_logic;                                        -- startofpacket
			src8_endofpacket    : out std_logic;                                        -- endofpacket
			src9_ready          : in  std_logic                     := 'X';             -- ready
			src9_valid          : out std_logic;                                        -- valid
			src9_data           : out std_logic_vector(75 downto 0);                    -- data
			src9_channel        : out std_logic_vector(13 downto 0);                    -- channel
			src9_startofpacket  : out std_logic;                                        -- startofpacket
			src9_endofpacket    : out std_logic;                                        -- endofpacket
			src10_ready         : in  std_logic                     := 'X';             -- ready
			src10_valid         : out std_logic;                                        -- valid
			src10_data          : out std_logic_vector(75 downto 0);                    -- data
			src10_channel       : out std_logic_vector(13 downto 0);                    -- channel
			src10_startofpacket : out std_logic;                                        -- startofpacket
			src10_endofpacket   : out std_logic;                                        -- endofpacket
			src11_ready         : in  std_logic                     := 'X';             -- ready
			src11_valid         : out std_logic;                                        -- valid
			src11_data          : out std_logic_vector(75 downto 0);                    -- data
			src11_channel       : out std_logic_vector(13 downto 0);                    -- channel
			src11_startofpacket : out std_logic;                                        -- startofpacket
			src11_endofpacket   : out std_logic;                                        -- endofpacket
			src12_ready         : in  std_logic                     := 'X';             -- ready
			src12_valid         : out std_logic;                                        -- valid
			src12_data          : out std_logic_vector(75 downto 0);                    -- data
			src12_channel       : out std_logic_vector(13 downto 0);                    -- channel
			src12_startofpacket : out std_logic;                                        -- startofpacket
			src12_endofpacket   : out std_logic;                                        -- endofpacket
			src13_ready         : in  std_logic                     := 'X';             -- ready
			src13_valid         : out std_logic;                                        -- valid
			src13_data          : out std_logic_vector(75 downto 0);                    -- data
			src13_channel       : out std_logic_vector(13 downto 0);                    -- channel
			src13_startofpacket : out std_logic;                                        -- startofpacket
			src13_endofpacket   : out std_logic                                         -- endofpacket
		);
	end component Nios1_cmd_xbar_demux_001;

	component Nios1_cmd_xbar_mux is
		port (
			clk                 : in  std_logic                     := 'X';             -- clk
			reset               : in  std_logic                     := 'X';             -- reset
			src_ready           : in  std_logic                     := 'X';             -- ready
			src_valid           : out std_logic;                                        -- valid
			src_data            : out std_logic_vector(75 downto 0);                    -- data
			src_channel         : out std_logic_vector(13 downto 0);                    -- channel
			src_startofpacket   : out std_logic;                                        -- startofpacket
			src_endofpacket     : out std_logic;                                        -- endofpacket
			sink0_ready         : out std_logic;                                        -- ready
			sink0_valid         : in  std_logic                     := 'X';             -- valid
			sink0_channel       : in  std_logic_vector(13 downto 0) := (others => 'X'); -- channel
			sink0_data          : in  std_logic_vector(75 downto 0) := (others => 'X'); -- data
			sink0_startofpacket : in  std_logic                     := 'X';             -- startofpacket
			sink0_endofpacket   : in  std_logic                     := 'X';             -- endofpacket
			sink1_ready         : out std_logic;                                        -- ready
			sink1_valid         : in  std_logic                     := 'X';             -- valid
			sink1_channel       : in  std_logic_vector(13 downto 0) := (others => 'X'); -- channel
			sink1_data          : in  std_logic_vector(75 downto 0) := (others => 'X'); -- data
			sink1_startofpacket : in  std_logic                     := 'X';             -- startofpacket
			sink1_endofpacket   : in  std_logic                     := 'X'              -- endofpacket
		);
	end component Nios1_cmd_xbar_mux;

	component Nios1_rsp_xbar_demux is
		port (
			clk                : in  std_logic                     := 'X';             -- clk
			reset              : in  std_logic                     := 'X';             -- reset
			sink_ready         : out std_logic;                                        -- ready
			sink_channel       : in  std_logic_vector(13 downto 0) := (others => 'X'); -- channel
			sink_data          : in  std_logic_vector(75 downto 0) := (others => 'X'); -- data
			sink_startofpacket : in  std_logic                     := 'X';             -- startofpacket
			sink_endofpacket   : in  std_logic                     := 'X';             -- endofpacket
			sink_valid         : in  std_logic_vector(0 downto 0)  := (others => 'X'); -- valid
			src0_ready         : in  std_logic                     := 'X';             -- ready
			src0_valid         : out std_logic;                                        -- valid
			src0_data          : out std_logic_vector(75 downto 0);                    -- data
			src0_channel       : out std_logic_vector(13 downto 0);                    -- channel
			src0_startofpacket : out std_logic;                                        -- startofpacket
			src0_endofpacket   : out std_logic;                                        -- endofpacket
			src1_ready         : in  std_logic                     := 'X';             -- ready
			src1_valid         : out std_logic;                                        -- valid
			src1_data          : out std_logic_vector(75 downto 0);                    -- data
			src1_channel       : out std_logic_vector(13 downto 0);                    -- channel
			src1_startofpacket : out std_logic;                                        -- startofpacket
			src1_endofpacket   : out std_logic                                         -- endofpacket
		);
	end component Nios1_rsp_xbar_demux;

	component Nios1_rsp_xbar_demux_002 is
		port (
			clk                : in  std_logic                     := 'X';             -- clk
			reset              : in  std_logic                     := 'X';             -- reset
			sink_ready         : out std_logic;                                        -- ready
			sink_channel       : in  std_logic_vector(13 downto 0) := (others => 'X'); -- channel
			sink_data          : in  std_logic_vector(75 downto 0) := (others => 'X'); -- data
			sink_startofpacket : in  std_logic                     := 'X';             -- startofpacket
			sink_endofpacket   : in  std_logic                     := 'X';             -- endofpacket
			sink_valid         : in  std_logic_vector(0 downto 0)  := (others => 'X'); -- valid
			src0_ready         : in  std_logic                     := 'X';             -- ready
			src0_valid         : out std_logic;                                        -- valid
			src0_data          : out std_logic_vector(75 downto 0);                    -- data
			src0_channel       : out std_logic_vector(13 downto 0);                    -- channel
			src0_startofpacket : out std_logic;                                        -- startofpacket
			src0_endofpacket   : out std_logic                                         -- endofpacket
		);
	end component Nios1_rsp_xbar_demux_002;

	component Nios1_rsp_xbar_mux is
		port (
			clk                 : in  std_logic                     := 'X';             -- clk
			reset               : in  std_logic                     := 'X';             -- reset
			src_ready           : in  std_logic                     := 'X';             -- ready
			src_valid           : out std_logic;                                        -- valid
			src_data            : out std_logic_vector(75 downto 0);                    -- data
			src_channel         : out std_logic_vector(13 downto 0);                    -- channel
			src_startofpacket   : out std_logic;                                        -- startofpacket
			src_endofpacket     : out std_logic;                                        -- endofpacket
			sink0_ready         : out std_logic;                                        -- ready
			sink0_valid         : in  std_logic                     := 'X';             -- valid
			sink0_channel       : in  std_logic_vector(13 downto 0) := (others => 'X'); -- channel
			sink0_data          : in  std_logic_vector(75 downto 0) := (others => 'X'); -- data
			sink0_startofpacket : in  std_logic                     := 'X';             -- startofpacket
			sink0_endofpacket   : in  std_logic                     := 'X';             -- endofpacket
			sink1_ready         : out std_logic;                                        -- ready
			sink1_valid         : in  std_logic                     := 'X';             -- valid
			sink1_channel       : in  std_logic_vector(13 downto 0) := (others => 'X'); -- channel
			sink1_data          : in  std_logic_vector(75 downto 0) := (others => 'X'); -- data
			sink1_startofpacket : in  std_logic                     := 'X';             -- startofpacket
			sink1_endofpacket   : in  std_logic                     := 'X'              -- endofpacket
		);
	end component Nios1_rsp_xbar_mux;

	component Nios1_rsp_xbar_mux_001 is
		port (
			clk                  : in  std_logic                     := 'X';             -- clk
			reset                : in  std_logic                     := 'X';             -- reset
			src_ready            : in  std_logic                     := 'X';             -- ready
			src_valid            : out std_logic;                                        -- valid
			src_data             : out std_logic_vector(75 downto 0);                    -- data
			src_channel          : out std_logic_vector(13 downto 0);                    -- channel
			src_startofpacket    : out std_logic;                                        -- startofpacket
			src_endofpacket      : out std_logic;                                        -- endofpacket
			sink0_ready          : out std_logic;                                        -- ready
			sink0_valid          : in  std_logic                     := 'X';             -- valid
			sink0_channel        : in  std_logic_vector(13 downto 0) := (others => 'X'); -- channel
			sink0_data           : in  std_logic_vector(75 downto 0) := (others => 'X'); -- data
			sink0_startofpacket  : in  std_logic                     := 'X';             -- startofpacket
			sink0_endofpacket    : in  std_logic                     := 'X';             -- endofpacket
			sink1_ready          : out std_logic;                                        -- ready
			sink1_valid          : in  std_logic                     := 'X';             -- valid
			sink1_channel        : in  std_logic_vector(13 downto 0) := (others => 'X'); -- channel
			sink1_data           : in  std_logic_vector(75 downto 0) := (others => 'X'); -- data
			sink1_startofpacket  : in  std_logic                     := 'X';             -- startofpacket
			sink1_endofpacket    : in  std_logic                     := 'X';             -- endofpacket
			sink2_ready          : out std_logic;                                        -- ready
			sink2_valid          : in  std_logic                     := 'X';             -- valid
			sink2_channel        : in  std_logic_vector(13 downto 0) := (others => 'X'); -- channel
			sink2_data           : in  std_logic_vector(75 downto 0) := (others => 'X'); -- data
			sink2_startofpacket  : in  std_logic                     := 'X';             -- startofpacket
			sink2_endofpacket    : in  std_logic                     := 'X';             -- endofpacket
			sink3_ready          : out std_logic;                                        -- ready
			sink3_valid          : in  std_logic                     := 'X';             -- valid
			sink3_channel        : in  std_logic_vector(13 downto 0) := (others => 'X'); -- channel
			sink3_data           : in  std_logic_vector(75 downto 0) := (others => 'X'); -- data
			sink3_startofpacket  : in  std_logic                     := 'X';             -- startofpacket
			sink3_endofpacket    : in  std_logic                     := 'X';             -- endofpacket
			sink4_ready          : out std_logic;                                        -- ready
			sink4_valid          : in  std_logic                     := 'X';             -- valid
			sink4_channel        : in  std_logic_vector(13 downto 0) := (others => 'X'); -- channel
			sink4_data           : in  std_logic_vector(75 downto 0) := (others => 'X'); -- data
			sink4_startofpacket  : in  std_logic                     := 'X';             -- startofpacket
			sink4_endofpacket    : in  std_logic                     := 'X';             -- endofpacket
			sink5_ready          : out std_logic;                                        -- ready
			sink5_valid          : in  std_logic                     := 'X';             -- valid
			sink5_channel        : in  std_logic_vector(13 downto 0) := (others => 'X'); -- channel
			sink5_data           : in  std_logic_vector(75 downto 0) := (others => 'X'); -- data
			sink5_startofpacket  : in  std_logic                     := 'X';             -- startofpacket
			sink5_endofpacket    : in  std_logic                     := 'X';             -- endofpacket
			sink6_ready          : out std_logic;                                        -- ready
			sink6_valid          : in  std_logic                     := 'X';             -- valid
			sink6_channel        : in  std_logic_vector(13 downto 0) := (others => 'X'); -- channel
			sink6_data           : in  std_logic_vector(75 downto 0) := (others => 'X'); -- data
			sink6_startofpacket  : in  std_logic                     := 'X';             -- startofpacket
			sink6_endofpacket    : in  std_logic                     := 'X';             -- endofpacket
			sink7_ready          : out std_logic;                                        -- ready
			sink7_valid          : in  std_logic                     := 'X';             -- valid
			sink7_channel        : in  std_logic_vector(13 downto 0) := (others => 'X'); -- channel
			sink7_data           : in  std_logic_vector(75 downto 0) := (others => 'X'); -- data
			sink7_startofpacket  : in  std_logic                     := 'X';             -- startofpacket
			sink7_endofpacket    : in  std_logic                     := 'X';             -- endofpacket
			sink8_ready          : out std_logic;                                        -- ready
			sink8_valid          : in  std_logic                     := 'X';             -- valid
			sink8_channel        : in  std_logic_vector(13 downto 0) := (others => 'X'); -- channel
			sink8_data           : in  std_logic_vector(75 downto 0) := (others => 'X'); -- data
			sink8_startofpacket  : in  std_logic                     := 'X';             -- startofpacket
			sink8_endofpacket    : in  std_logic                     := 'X';             -- endofpacket
			sink9_ready          : out std_logic;                                        -- ready
			sink9_valid          : in  std_logic                     := 'X';             -- valid
			sink9_channel        : in  std_logic_vector(13 downto 0) := (others => 'X'); -- channel
			sink9_data           : in  std_logic_vector(75 downto 0) := (others => 'X'); -- data
			sink9_startofpacket  : in  std_logic                     := 'X';             -- startofpacket
			sink9_endofpacket    : in  std_logic                     := 'X';             -- endofpacket
			sink10_ready         : out std_logic;                                        -- ready
			sink10_valid         : in  std_logic                     := 'X';             -- valid
			sink10_channel       : in  std_logic_vector(13 downto 0) := (others => 'X'); -- channel
			sink10_data          : in  std_logic_vector(75 downto 0) := (others => 'X'); -- data
			sink10_startofpacket : in  std_logic                     := 'X';             -- startofpacket
			sink10_endofpacket   : in  std_logic                     := 'X';             -- endofpacket
			sink11_ready         : out std_logic;                                        -- ready
			sink11_valid         : in  std_logic                     := 'X';             -- valid
			sink11_channel       : in  std_logic_vector(13 downto 0) := (others => 'X'); -- channel
			sink11_data          : in  std_logic_vector(75 downto 0) := (others => 'X'); -- data
			sink11_startofpacket : in  std_logic                     := 'X';             -- startofpacket
			sink11_endofpacket   : in  std_logic                     := 'X';             -- endofpacket
			sink12_ready         : out std_logic;                                        -- ready
			sink12_valid         : in  std_logic                     := 'X';             -- valid
			sink12_channel       : in  std_logic_vector(13 downto 0) := (others => 'X'); -- channel
			sink12_data          : in  std_logic_vector(75 downto 0) := (others => 'X'); -- data
			sink12_startofpacket : in  std_logic                     := 'X';             -- startofpacket
			sink12_endofpacket   : in  std_logic                     := 'X';             -- endofpacket
			sink13_ready         : out std_logic;                                        -- ready
			sink13_valid         : in  std_logic                     := 'X';             -- valid
			sink13_channel       : in  std_logic_vector(13 downto 0) := (others => 'X'); -- channel
			sink13_data          : in  std_logic_vector(75 downto 0) := (others => 'X'); -- data
			sink13_startofpacket : in  std_logic                     := 'X';             -- startofpacket
			sink13_endofpacket   : in  std_logic                     := 'X'              -- endofpacket
		);
	end component Nios1_rsp_xbar_mux_001;

	component Nios1_irq_mapper is
		port (
			clk           : in  std_logic                     := 'X'; -- clk
			reset         : in  std_logic                     := 'X'; -- reset
			receiver0_irq : in  std_logic                     := 'X'; -- irq
			receiver1_irq : in  std_logic                     := 'X'; -- irq
			receiver2_irq : in  std_logic                     := 'X'; -- irq
			receiver3_irq : in  std_logic                     := 'X'; -- irq
			receiver4_irq : in  std_logic                     := 'X'; -- irq
			sender_irq    : out std_logic_vector(31 downto 0)         -- irq
		);
	end component Nios1_irq_mapper;

	signal nios2_qsys_instruction_master_waitrequest                                                         : std_logic;                     -- nios2_qsys_instruction_master_translator:av_waitrequest -> nios2_qsys:i_waitrequest
	signal nios2_qsys_instruction_master_address                                                             : std_logic_vector(18 downto 0); -- nios2_qsys:i_address -> nios2_qsys_instruction_master_translator:av_address
	signal nios2_qsys_instruction_master_read                                                                : std_logic;                     -- nios2_qsys:i_read -> nios2_qsys_instruction_master_translator:av_read
	signal nios2_qsys_instruction_master_readdata                                                            : std_logic_vector(31 downto 0); -- nios2_qsys_instruction_master_translator:av_readdata -> nios2_qsys:i_readdata
	signal nios2_qsys_instruction_master_readdatavalid                                                       : std_logic;                     -- nios2_qsys_instruction_master_translator:av_readdatavalid -> nios2_qsys:i_readdatavalid
	signal nios2_qsys_data_master_waitrequest                                                                : std_logic;                     -- nios2_qsys_data_master_translator:av_waitrequest -> nios2_qsys:d_waitrequest
	signal nios2_qsys_data_master_writedata                                                                  : std_logic_vector(31 downto 0); -- nios2_qsys:d_writedata -> nios2_qsys_data_master_translator:av_writedata
	signal nios2_qsys_data_master_address                                                                    : std_logic_vector(18 downto 0); -- nios2_qsys:d_address -> nios2_qsys_data_master_translator:av_address
	signal nios2_qsys_data_master_write                                                                      : std_logic;                     -- nios2_qsys:d_write -> nios2_qsys_data_master_translator:av_write
	signal nios2_qsys_data_master_read                                                                       : std_logic;                     -- nios2_qsys:d_read -> nios2_qsys_data_master_translator:av_read
	signal nios2_qsys_data_master_readdata                                                                   : std_logic_vector(31 downto 0); -- nios2_qsys_data_master_translator:av_readdata -> nios2_qsys:d_readdata
	signal nios2_qsys_data_master_debugaccess                                                                : std_logic;                     -- nios2_qsys:jtag_debug_module_debugaccess_to_roms -> nios2_qsys_data_master_translator:av_debugaccess
	signal nios2_qsys_data_master_readdatavalid                                                              : std_logic;                     -- nios2_qsys_data_master_translator:av_readdatavalid -> nios2_qsys:d_readdatavalid
	signal nios2_qsys_data_master_byteenable                                                                 : std_logic_vector(3 downto 0);  -- nios2_qsys:d_byteenable -> nios2_qsys_data_master_translator:av_byteenable
	signal nios2_qsys_jtag_debug_module_translator_avalon_anti_slave_0_writedata                             : std_logic_vector(31 downto 0); -- nios2_qsys_jtag_debug_module_translator:av_writedata -> nios2_qsys:jtag_debug_module_writedata
	signal nios2_qsys_jtag_debug_module_translator_avalon_anti_slave_0_address                               : std_logic_vector(8 downto 0);  -- nios2_qsys_jtag_debug_module_translator:av_address -> nios2_qsys:jtag_debug_module_address
	signal nios2_qsys_jtag_debug_module_translator_avalon_anti_slave_0_chipselect                            : std_logic;                     -- nios2_qsys_jtag_debug_module_translator:av_chipselect -> nios2_qsys:jtag_debug_module_select
	signal nios2_qsys_jtag_debug_module_translator_avalon_anti_slave_0_write                                 : std_logic;                     -- nios2_qsys_jtag_debug_module_translator:av_write -> nios2_qsys:jtag_debug_module_write
	signal nios2_qsys_jtag_debug_module_translator_avalon_anti_slave_0_readdata                              : std_logic_vector(31 downto 0); -- nios2_qsys:jtag_debug_module_readdata -> nios2_qsys_jtag_debug_module_translator:av_readdata
	signal nios2_qsys_jtag_debug_module_translator_avalon_anti_slave_0_begintransfer                         : std_logic;                     -- nios2_qsys_jtag_debug_module_translator:av_begintransfer -> nios2_qsys:jtag_debug_module_begintransfer
	signal nios2_qsys_jtag_debug_module_translator_avalon_anti_slave_0_debugaccess                           : std_logic;                     -- nios2_qsys_jtag_debug_module_translator:av_debugaccess -> nios2_qsys:jtag_debug_module_debugaccess
	signal nios2_qsys_jtag_debug_module_translator_avalon_anti_slave_0_byteenable                            : std_logic_vector(3 downto 0);  -- nios2_qsys_jtag_debug_module_translator:av_byteenable -> nios2_qsys:jtag_debug_module_byteenable
	signal onchip_memory_s1_translator_avalon_anti_slave_0_writedata                                         : std_logic_vector(31 downto 0); -- onchip_memory_s1_translator:av_writedata -> onchip_memory:writedata
	signal onchip_memory_s1_translator_avalon_anti_slave_0_address                                           : std_logic_vector(14 downto 0); -- onchip_memory_s1_translator:av_address -> onchip_memory:address
	signal onchip_memory_s1_translator_avalon_anti_slave_0_chipselect                                        : std_logic;                     -- onchip_memory_s1_translator:av_chipselect -> onchip_memory:chipselect
	signal onchip_memory_s1_translator_avalon_anti_slave_0_clken                                             : std_logic;                     -- onchip_memory_s1_translator:av_clken -> onchip_memory:clken
	signal onchip_memory_s1_translator_avalon_anti_slave_0_write                                             : std_logic;                     -- onchip_memory_s1_translator:av_write -> onchip_memory:write
	signal onchip_memory_s1_translator_avalon_anti_slave_0_readdata                                          : std_logic_vector(31 downto 0); -- onchip_memory:readdata -> onchip_memory_s1_translator:av_readdata
	signal onchip_memory_s1_translator_avalon_anti_slave_0_byteenable                                        : std_logic_vector(3 downto 0);  -- onchip_memory_s1_translator:av_byteenable -> onchip_memory:byteenable
	signal jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_waitrequest                            : std_logic;                     -- jtag_uart:av_waitrequest -> jtag_uart_avalon_jtag_slave_translator:av_waitrequest
	signal jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_writedata                              : std_logic_vector(31 downto 0); -- jtag_uart_avalon_jtag_slave_translator:av_writedata -> jtag_uart:av_writedata
	signal jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_address                                : std_logic;                     -- jtag_uart_avalon_jtag_slave_translator:av_address -> jtag_uart:av_address
	signal jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_chipselect                             : std_logic;                     -- jtag_uart_avalon_jtag_slave_translator:av_chipselect -> jtag_uart:av_chipselect
	signal jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_write                                  : std_logic;                     -- jtag_uart_avalon_jtag_slave_translator:av_write -> jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_write:in
	signal jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_read                                   : std_logic;                     -- jtag_uart_avalon_jtag_slave_translator:av_read -> jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_read:in
	signal jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_readdata                               : std_logic_vector(31 downto 0); -- jtag_uart:av_readdata -> jtag_uart_avalon_jtag_slave_translator:av_readdata
	signal sysid_qsys_control_slave_translator_avalon_anti_slave_0_address                                   : std_logic;                     -- sysid_qsys_control_slave_translator:av_address -> sysid_qsys:address
	signal sysid_qsys_control_slave_translator_avalon_anti_slave_0_readdata                                  : std_logic_vector(31 downto 0); -- sysid_qsys:readdata -> sysid_qsys_control_slave_translator:av_readdata
	signal pio_ledg_s1_translator_avalon_anti_slave_0_writedata                                              : std_logic_vector(31 downto 0); -- pio_LEDG_s1_translator:av_writedata -> pio_LEDG:writedata
	signal pio_ledg_s1_translator_avalon_anti_slave_0_address                                                : std_logic_vector(2 downto 0);  -- pio_LEDG_s1_translator:av_address -> pio_LEDG:address
	signal pio_ledg_s1_translator_avalon_anti_slave_0_chipselect                                             : std_logic;                     -- pio_LEDG_s1_translator:av_chipselect -> pio_LEDG:chipselect
	signal pio_ledg_s1_translator_avalon_anti_slave_0_write                                                  : std_logic;                     -- pio_LEDG_s1_translator:av_write -> pio_ledg_s1_translator_avalon_anti_slave_0_write:in
	signal pio_ledg_s1_translator_avalon_anti_slave_0_readdata                                               : std_logic_vector(31 downto 0); -- pio_LEDG:readdata -> pio_LEDG_s1_translator:av_readdata
	signal pio_ledr_s1_translator_avalon_anti_slave_0_writedata                                              : std_logic_vector(31 downto 0); -- pio_LEDR_s1_translator:av_writedata -> pio_LEDR:writedata
	signal pio_ledr_s1_translator_avalon_anti_slave_0_address                                                : std_logic_vector(2 downto 0);  -- pio_LEDR_s1_translator:av_address -> pio_LEDR:address
	signal pio_ledr_s1_translator_avalon_anti_slave_0_chipselect                                             : std_logic;                     -- pio_LEDR_s1_translator:av_chipselect -> pio_LEDR:chipselect
	signal pio_ledr_s1_translator_avalon_anti_slave_0_write                                                  : std_logic;                     -- pio_LEDR_s1_translator:av_write -> pio_ledr_s1_translator_avalon_anti_slave_0_write:in
	signal pio_ledr_s1_translator_avalon_anti_slave_0_readdata                                               : std_logic_vector(31 downto 0); -- pio_LEDR:readdata -> pio_LEDR_s1_translator:av_readdata
	signal pio_sw_s1_translator_avalon_anti_slave_0_address                                                  : std_logic_vector(1 downto 0);  -- pio_SW_s1_translator:av_address -> pio_SW:address
	signal pio_sw_s1_translator_avalon_anti_slave_0_readdata                                                 : std_logic_vector(31 downto 0); -- pio_SW:readdata -> pio_SW_s1_translator:av_readdata
	signal pio_button_s1_translator_avalon_anti_slave_0_writedata                                            : std_logic_vector(31 downto 0); -- pio_Button_s1_translator:av_writedata -> pio_Button:writedata
	signal pio_button_s1_translator_avalon_anti_slave_0_address                                              : std_logic_vector(1 downto 0);  -- pio_Button_s1_translator:av_address -> pio_Button:address
	signal pio_button_s1_translator_avalon_anti_slave_0_chipselect                                           : std_logic;                     -- pio_Button_s1_translator:av_chipselect -> pio_Button:chipselect
	signal pio_button_s1_translator_avalon_anti_slave_0_write                                                : std_logic;                     -- pio_Button_s1_translator:av_write -> pio_button_s1_translator_avalon_anti_slave_0_write:in
	signal pio_button_s1_translator_avalon_anti_slave_0_readdata                                             : std_logic_vector(31 downto 0); -- pio_Button:readdata -> pio_Button_s1_translator:av_readdata
	signal lcd_control_slave_translator_avalon_anti_slave_0_writedata                                        : std_logic_vector(7 downto 0);  -- lcd_control_slave_translator:av_writedata -> lcd:writedata
	signal lcd_control_slave_translator_avalon_anti_slave_0_address                                          : std_logic_vector(1 downto 0);  -- lcd_control_slave_translator:av_address -> lcd:address
	signal lcd_control_slave_translator_avalon_anti_slave_0_write                                            : std_logic;                     -- lcd_control_slave_translator:av_write -> lcd:write
	signal lcd_control_slave_translator_avalon_anti_slave_0_read                                             : std_logic;                     -- lcd_control_slave_translator:av_read -> lcd:read
	signal lcd_control_slave_translator_avalon_anti_slave_0_readdata                                         : std_logic_vector(7 downto 0);  -- lcd:readdata -> lcd_control_slave_translator:av_readdata
	signal lcd_control_slave_translator_avalon_anti_slave_0_begintransfer                                    : std_logic;                     -- lcd_control_slave_translator:av_begintransfer -> lcd:begintransfer
	signal uart_s1_translator_avalon_anti_slave_0_writedata                                                  : std_logic_vector(15 downto 0); -- uart_s1_translator:av_writedata -> uart:writedata
	signal uart_s1_translator_avalon_anti_slave_0_address                                                    : std_logic_vector(2 downto 0);  -- uart_s1_translator:av_address -> uart:address
	signal uart_s1_translator_avalon_anti_slave_0_chipselect                                                 : std_logic;                     -- uart_s1_translator:av_chipselect -> uart:chipselect
	signal uart_s1_translator_avalon_anti_slave_0_write                                                      : std_logic;                     -- uart_s1_translator:av_write -> uart_s1_translator_avalon_anti_slave_0_write:in
	signal uart_s1_translator_avalon_anti_slave_0_read                                                       : std_logic;                     -- uart_s1_translator:av_read -> uart_s1_translator_avalon_anti_slave_0_read:in
	signal uart_s1_translator_avalon_anti_slave_0_readdata                                                   : std_logic_vector(15 downto 0); -- uart:readdata -> uart_s1_translator:av_readdata
	signal uart_s1_translator_avalon_anti_slave_0_begintransfer                                              : std_logic;                     -- uart_s1_translator:av_begintransfer -> uart:begintransfer
	signal timer_0_s1_translator_avalon_anti_slave_0_writedata                                               : std_logic_vector(15 downto 0); -- timer_0_s1_translator:av_writedata -> timer_0:writedata
	signal timer_0_s1_translator_avalon_anti_slave_0_address                                                 : std_logic_vector(2 downto 0);  -- timer_0_s1_translator:av_address -> timer_0:address
	signal timer_0_s1_translator_avalon_anti_slave_0_chipselect                                              : std_logic;                     -- timer_0_s1_translator:av_chipselect -> timer_0:chipselect
	signal timer_0_s1_translator_avalon_anti_slave_0_write                                                   : std_logic;                     -- timer_0_s1_translator:av_write -> timer_0_s1_translator_avalon_anti_slave_0_write:in
	signal timer_0_s1_translator_avalon_anti_slave_0_readdata                                                : std_logic_vector(15 downto 0); -- timer_0:readdata -> timer_0_s1_translator:av_readdata
	signal pio_data_s1_translator_avalon_anti_slave_0_address                                                : std_logic_vector(1 downto 0);  -- pio_Data_s1_translator:av_address -> pio_Data:address
	signal pio_data_s1_translator_avalon_anti_slave_0_readdata                                               : std_logic_vector(31 downto 0); -- pio_Data:readdata -> pio_Data_s1_translator:av_readdata
	signal pio_rdydata_s1_translator_avalon_anti_slave_0_writedata                                           : std_logic_vector(31 downto 0); -- pio_RdyData_s1_translator:av_writedata -> pio_RdyData:writedata
	signal pio_rdydata_s1_translator_avalon_anti_slave_0_address                                             : std_logic_vector(1 downto 0);  -- pio_RdyData_s1_translator:av_address -> pio_RdyData:address
	signal pio_rdydata_s1_translator_avalon_anti_slave_0_chipselect                                          : std_logic;                     -- pio_RdyData_s1_translator:av_chipselect -> pio_RdyData:chipselect
	signal pio_rdydata_s1_translator_avalon_anti_slave_0_write                                               : std_logic;                     -- pio_RdyData_s1_translator:av_write -> pio_rdydata_s1_translator_avalon_anti_slave_0_write:in
	signal pio_rdydata_s1_translator_avalon_anti_slave_0_readdata                                            : std_logic_vector(31 downto 0); -- pio_RdyData:readdata -> pio_RdyData_s1_translator:av_readdata
	signal pio_dataread_s1_translator_avalon_anti_slave_0_writedata                                          : std_logic_vector(31 downto 0); -- pio_DataRead_s1_translator:av_writedata -> pio_DataRead:writedata
	signal pio_dataread_s1_translator_avalon_anti_slave_0_address                                            : std_logic_vector(2 downto 0);  -- pio_DataRead_s1_translator:av_address -> pio_DataRead:address
	signal pio_dataread_s1_translator_avalon_anti_slave_0_chipselect                                         : std_logic;                     -- pio_DataRead_s1_translator:av_chipselect -> pio_DataRead:chipselect
	signal pio_dataread_s1_translator_avalon_anti_slave_0_write                                              : std_logic;                     -- pio_DataRead_s1_translator:av_write -> pio_dataread_s1_translator_avalon_anti_slave_0_write:in
	signal pio_dataread_s1_translator_avalon_anti_slave_0_readdata                                           : std_logic_vector(31 downto 0); -- pio_DataRead:readdata -> pio_DataRead_s1_translator:av_readdata
	signal pio_ledg_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest                              : std_logic;                     -- pio_LEDG_s1_translator:uav_waitrequest -> pio_LEDG_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	signal pio_ledg_s1_translator_avalon_universal_slave_0_agent_m0_burstcount                               : std_logic_vector(2 downto 0);  -- pio_LEDG_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> pio_LEDG_s1_translator:uav_burstcount
	signal pio_ledg_s1_translator_avalon_universal_slave_0_agent_m0_writedata                                : std_logic_vector(31 downto 0); -- pio_LEDG_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> pio_LEDG_s1_translator:uav_writedata
	signal pio_ledg_s1_translator_avalon_universal_slave_0_agent_m0_address                                  : std_logic_vector(18 downto 0); -- pio_LEDG_s1_translator_avalon_universal_slave_0_agent:m0_address -> pio_LEDG_s1_translator:uav_address
	signal pio_ledg_s1_translator_avalon_universal_slave_0_agent_m0_write                                    : std_logic;                     -- pio_LEDG_s1_translator_avalon_universal_slave_0_agent:m0_write -> pio_LEDG_s1_translator:uav_write
	signal pio_ledg_s1_translator_avalon_universal_slave_0_agent_m0_lock                                     : std_logic;                     -- pio_LEDG_s1_translator_avalon_universal_slave_0_agent:m0_lock -> pio_LEDG_s1_translator:uav_lock
	signal pio_ledg_s1_translator_avalon_universal_slave_0_agent_m0_read                                     : std_logic;                     -- pio_LEDG_s1_translator_avalon_universal_slave_0_agent:m0_read -> pio_LEDG_s1_translator:uav_read
	signal pio_ledg_s1_translator_avalon_universal_slave_0_agent_m0_readdata                                 : std_logic_vector(31 downto 0); -- pio_LEDG_s1_translator:uav_readdata -> pio_LEDG_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	signal pio_ledg_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid                            : std_logic;                     -- pio_LEDG_s1_translator:uav_readdatavalid -> pio_LEDG_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	signal pio_ledg_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess                              : std_logic;                     -- pio_LEDG_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> pio_LEDG_s1_translator:uav_debugaccess
	signal pio_ledg_s1_translator_avalon_universal_slave_0_agent_m0_byteenable                               : std_logic_vector(3 downto 0);  -- pio_LEDG_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> pio_LEDG_s1_translator:uav_byteenable
	signal pio_ledg_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket                       : std_logic;                     -- pio_LEDG_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> pio_LEDG_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	signal pio_ledg_s1_translator_avalon_universal_slave_0_agent_rf_source_valid                             : std_logic;                     -- pio_LEDG_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> pio_LEDG_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	signal pio_ledg_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket                     : std_logic;                     -- pio_LEDG_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> pio_LEDG_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	signal pio_ledg_s1_translator_avalon_universal_slave_0_agent_rf_source_data                              : std_logic_vector(76 downto 0); -- pio_LEDG_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> pio_LEDG_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	signal pio_ledg_s1_translator_avalon_universal_slave_0_agent_rf_source_ready                             : std_logic;                     -- pio_LEDG_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> pio_LEDG_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	signal pio_ledg_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket                    : std_logic;                     -- pio_LEDG_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> pio_LEDG_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	signal pio_ledg_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid                          : std_logic;                     -- pio_LEDG_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> pio_LEDG_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	signal pio_ledg_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket                  : std_logic;                     -- pio_LEDG_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> pio_LEDG_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	signal pio_ledg_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data                           : std_logic_vector(76 downto 0); -- pio_LEDG_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> pio_LEDG_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	signal pio_ledg_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready                          : std_logic;                     -- pio_LEDG_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> pio_LEDG_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	signal pio_ledg_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid                        : std_logic;                     -- pio_LEDG_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> pio_LEDG_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	signal pio_ledg_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data                         : std_logic_vector(31 downto 0); -- pio_LEDG_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> pio_LEDG_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	signal pio_ledg_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready                        : std_logic;                     -- pio_LEDG_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> pio_LEDG_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	signal pio_ledr_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest                              : std_logic;                     -- pio_LEDR_s1_translator:uav_waitrequest -> pio_LEDR_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	signal pio_ledr_s1_translator_avalon_universal_slave_0_agent_m0_burstcount                               : std_logic_vector(2 downto 0);  -- pio_LEDR_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> pio_LEDR_s1_translator:uav_burstcount
	signal pio_ledr_s1_translator_avalon_universal_slave_0_agent_m0_writedata                                : std_logic_vector(31 downto 0); -- pio_LEDR_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> pio_LEDR_s1_translator:uav_writedata
	signal pio_ledr_s1_translator_avalon_universal_slave_0_agent_m0_address                                  : std_logic_vector(18 downto 0); -- pio_LEDR_s1_translator_avalon_universal_slave_0_agent:m0_address -> pio_LEDR_s1_translator:uav_address
	signal pio_ledr_s1_translator_avalon_universal_slave_0_agent_m0_write                                    : std_logic;                     -- pio_LEDR_s1_translator_avalon_universal_slave_0_agent:m0_write -> pio_LEDR_s1_translator:uav_write
	signal pio_ledr_s1_translator_avalon_universal_slave_0_agent_m0_lock                                     : std_logic;                     -- pio_LEDR_s1_translator_avalon_universal_slave_0_agent:m0_lock -> pio_LEDR_s1_translator:uav_lock
	signal pio_ledr_s1_translator_avalon_universal_slave_0_agent_m0_read                                     : std_logic;                     -- pio_LEDR_s1_translator_avalon_universal_slave_0_agent:m0_read -> pio_LEDR_s1_translator:uav_read
	signal pio_ledr_s1_translator_avalon_universal_slave_0_agent_m0_readdata                                 : std_logic_vector(31 downto 0); -- pio_LEDR_s1_translator:uav_readdata -> pio_LEDR_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	signal pio_ledr_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid                            : std_logic;                     -- pio_LEDR_s1_translator:uav_readdatavalid -> pio_LEDR_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	signal pio_ledr_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess                              : std_logic;                     -- pio_LEDR_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> pio_LEDR_s1_translator:uav_debugaccess
	signal pio_ledr_s1_translator_avalon_universal_slave_0_agent_m0_byteenable                               : std_logic_vector(3 downto 0);  -- pio_LEDR_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> pio_LEDR_s1_translator:uav_byteenable
	signal pio_ledr_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket                       : std_logic;                     -- pio_LEDR_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> pio_LEDR_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	signal pio_ledr_s1_translator_avalon_universal_slave_0_agent_rf_source_valid                             : std_logic;                     -- pio_LEDR_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> pio_LEDR_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	signal pio_ledr_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket                     : std_logic;                     -- pio_LEDR_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> pio_LEDR_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	signal pio_ledr_s1_translator_avalon_universal_slave_0_agent_rf_source_data                              : std_logic_vector(76 downto 0); -- pio_LEDR_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> pio_LEDR_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	signal pio_ledr_s1_translator_avalon_universal_slave_0_agent_rf_source_ready                             : std_logic;                     -- pio_LEDR_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> pio_LEDR_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	signal pio_ledr_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket                    : std_logic;                     -- pio_LEDR_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> pio_LEDR_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	signal pio_ledr_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid                          : std_logic;                     -- pio_LEDR_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> pio_LEDR_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	signal pio_ledr_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket                  : std_logic;                     -- pio_LEDR_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> pio_LEDR_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	signal pio_ledr_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data                           : std_logic_vector(76 downto 0); -- pio_LEDR_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> pio_LEDR_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	signal pio_ledr_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready                          : std_logic;                     -- pio_LEDR_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> pio_LEDR_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	signal pio_ledr_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid                        : std_logic;                     -- pio_LEDR_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> pio_LEDR_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	signal pio_ledr_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data                         : std_logic_vector(31 downto 0); -- pio_LEDR_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> pio_LEDR_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	signal pio_ledr_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready                        : std_logic;                     -- pio_LEDR_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> pio_LEDR_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	signal sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest                 : std_logic;                     -- sysid_qsys_control_slave_translator:uav_waitrequest -> sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent:m0_waitrequest
	signal sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent_m0_burstcount                  : std_logic_vector(2 downto 0);  -- sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent:m0_burstcount -> sysid_qsys_control_slave_translator:uav_burstcount
	signal sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent_m0_writedata                   : std_logic_vector(31 downto 0); -- sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent:m0_writedata -> sysid_qsys_control_slave_translator:uav_writedata
	signal sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent_m0_address                     : std_logic_vector(18 downto 0); -- sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent:m0_address -> sysid_qsys_control_slave_translator:uav_address
	signal sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent_m0_write                       : std_logic;                     -- sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent:m0_write -> sysid_qsys_control_slave_translator:uav_write
	signal sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent_m0_lock                        : std_logic;                     -- sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent:m0_lock -> sysid_qsys_control_slave_translator:uav_lock
	signal sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent_m0_read                        : std_logic;                     -- sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent:m0_read -> sysid_qsys_control_slave_translator:uav_read
	signal sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent_m0_readdata                    : std_logic_vector(31 downto 0); -- sysid_qsys_control_slave_translator:uav_readdata -> sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent:m0_readdata
	signal sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid               : std_logic;                     -- sysid_qsys_control_slave_translator:uav_readdatavalid -> sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	signal sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess                 : std_logic;                     -- sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent:m0_debugaccess -> sysid_qsys_control_slave_translator:uav_debugaccess
	signal sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent_m0_byteenable                  : std_logic_vector(3 downto 0);  -- sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent:m0_byteenable -> sysid_qsys_control_slave_translator:uav_byteenable
	signal sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket          : std_logic;                     -- sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	signal sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent_rf_source_valid                : std_logic;                     -- sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent:rf_source_valid -> sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	signal sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket        : std_logic;                     -- sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	signal sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent_rf_source_data                 : std_logic_vector(76 downto 0); -- sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent:rf_source_data -> sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	signal sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent_rf_source_ready                : std_logic;                     -- sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent:rf_source_ready
	signal sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket       : std_logic;                     -- sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	signal sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid             : std_logic;                     -- sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent:rf_sink_valid
	signal sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket     : std_logic;                     -- sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	signal sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data              : std_logic_vector(76 downto 0); -- sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent:rf_sink_data
	signal sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready             : std_logic;                     -- sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent:rf_sink_ready -> sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	signal sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid           : std_logic;                     -- sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	signal sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data            : std_logic_vector(31 downto 0); -- sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	signal sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready           : std_logic;                     -- sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	signal pio_dataread_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest                          : std_logic;                     -- pio_DataRead_s1_translator:uav_waitrequest -> pio_DataRead_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	signal pio_dataread_s1_translator_avalon_universal_slave_0_agent_m0_burstcount                           : std_logic_vector(2 downto 0);  -- pio_DataRead_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> pio_DataRead_s1_translator:uav_burstcount
	signal pio_dataread_s1_translator_avalon_universal_slave_0_agent_m0_writedata                            : std_logic_vector(31 downto 0); -- pio_DataRead_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> pio_DataRead_s1_translator:uav_writedata
	signal pio_dataread_s1_translator_avalon_universal_slave_0_agent_m0_address                              : std_logic_vector(18 downto 0); -- pio_DataRead_s1_translator_avalon_universal_slave_0_agent:m0_address -> pio_DataRead_s1_translator:uav_address
	signal pio_dataread_s1_translator_avalon_universal_slave_0_agent_m0_write                                : std_logic;                     -- pio_DataRead_s1_translator_avalon_universal_slave_0_agent:m0_write -> pio_DataRead_s1_translator:uav_write
	signal pio_dataread_s1_translator_avalon_universal_slave_0_agent_m0_lock                                 : std_logic;                     -- pio_DataRead_s1_translator_avalon_universal_slave_0_agent:m0_lock -> pio_DataRead_s1_translator:uav_lock
	signal pio_dataread_s1_translator_avalon_universal_slave_0_agent_m0_read                                 : std_logic;                     -- pio_DataRead_s1_translator_avalon_universal_slave_0_agent:m0_read -> pio_DataRead_s1_translator:uav_read
	signal pio_dataread_s1_translator_avalon_universal_slave_0_agent_m0_readdata                             : std_logic_vector(31 downto 0); -- pio_DataRead_s1_translator:uav_readdata -> pio_DataRead_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	signal pio_dataread_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid                        : std_logic;                     -- pio_DataRead_s1_translator:uav_readdatavalid -> pio_DataRead_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	signal pio_dataread_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess                          : std_logic;                     -- pio_DataRead_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> pio_DataRead_s1_translator:uav_debugaccess
	signal pio_dataread_s1_translator_avalon_universal_slave_0_agent_m0_byteenable                           : std_logic_vector(3 downto 0);  -- pio_DataRead_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> pio_DataRead_s1_translator:uav_byteenable
	signal pio_dataread_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket                   : std_logic;                     -- pio_DataRead_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> pio_DataRead_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	signal pio_dataread_s1_translator_avalon_universal_slave_0_agent_rf_source_valid                         : std_logic;                     -- pio_DataRead_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> pio_DataRead_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	signal pio_dataread_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket                 : std_logic;                     -- pio_DataRead_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> pio_DataRead_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	signal pio_dataread_s1_translator_avalon_universal_slave_0_agent_rf_source_data                          : std_logic_vector(76 downto 0); -- pio_DataRead_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> pio_DataRead_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	signal pio_dataread_s1_translator_avalon_universal_slave_0_agent_rf_source_ready                         : std_logic;                     -- pio_DataRead_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> pio_DataRead_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	signal pio_dataread_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket                : std_logic;                     -- pio_DataRead_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> pio_DataRead_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	signal pio_dataread_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid                      : std_logic;                     -- pio_DataRead_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> pio_DataRead_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	signal pio_dataread_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket              : std_logic;                     -- pio_DataRead_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> pio_DataRead_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	signal pio_dataread_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data                       : std_logic_vector(76 downto 0); -- pio_DataRead_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> pio_DataRead_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	signal pio_dataread_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready                      : std_logic;                     -- pio_DataRead_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> pio_DataRead_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	signal pio_dataread_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid                    : std_logic;                     -- pio_DataRead_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> pio_DataRead_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	signal pio_dataread_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data                     : std_logic_vector(31 downto 0); -- pio_DataRead_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> pio_DataRead_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	signal pio_dataread_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready                    : std_logic;                     -- pio_DataRead_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> pio_DataRead_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	signal nios2_qsys_data_master_translator_avalon_universal_master_0_waitrequest                           : std_logic;                     -- nios2_qsys_data_master_translator_avalon_universal_master_0_agent:av_waitrequest -> nios2_qsys_data_master_translator:uav_waitrequest
	signal nios2_qsys_data_master_translator_avalon_universal_master_0_burstcount                            : std_logic_vector(2 downto 0);  -- nios2_qsys_data_master_translator:uav_burstcount -> nios2_qsys_data_master_translator_avalon_universal_master_0_agent:av_burstcount
	signal nios2_qsys_data_master_translator_avalon_universal_master_0_writedata                             : std_logic_vector(31 downto 0); -- nios2_qsys_data_master_translator:uav_writedata -> nios2_qsys_data_master_translator_avalon_universal_master_0_agent:av_writedata
	signal nios2_qsys_data_master_translator_avalon_universal_master_0_address                               : std_logic_vector(18 downto 0); -- nios2_qsys_data_master_translator:uav_address -> nios2_qsys_data_master_translator_avalon_universal_master_0_agent:av_address
	signal nios2_qsys_data_master_translator_avalon_universal_master_0_lock                                  : std_logic;                     -- nios2_qsys_data_master_translator:uav_lock -> nios2_qsys_data_master_translator_avalon_universal_master_0_agent:av_lock
	signal nios2_qsys_data_master_translator_avalon_universal_master_0_write                                 : std_logic;                     -- nios2_qsys_data_master_translator:uav_write -> nios2_qsys_data_master_translator_avalon_universal_master_0_agent:av_write
	signal nios2_qsys_data_master_translator_avalon_universal_master_0_read                                  : std_logic;                     -- nios2_qsys_data_master_translator:uav_read -> nios2_qsys_data_master_translator_avalon_universal_master_0_agent:av_read
	signal nios2_qsys_data_master_translator_avalon_universal_master_0_readdata                              : std_logic_vector(31 downto 0); -- nios2_qsys_data_master_translator_avalon_universal_master_0_agent:av_readdata -> nios2_qsys_data_master_translator:uav_readdata
	signal nios2_qsys_data_master_translator_avalon_universal_master_0_debugaccess                           : std_logic;                     -- nios2_qsys_data_master_translator:uav_debugaccess -> nios2_qsys_data_master_translator_avalon_universal_master_0_agent:av_debugaccess
	signal nios2_qsys_data_master_translator_avalon_universal_master_0_byteenable                            : std_logic_vector(3 downto 0);  -- nios2_qsys_data_master_translator:uav_byteenable -> nios2_qsys_data_master_translator_avalon_universal_master_0_agent:av_byteenable
	signal nios2_qsys_data_master_translator_avalon_universal_master_0_readdatavalid                         : std_logic;                     -- nios2_qsys_data_master_translator_avalon_universal_master_0_agent:av_readdatavalid -> nios2_qsys_data_master_translator:uav_readdatavalid
	signal lcd_control_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest                        : std_logic;                     -- lcd_control_slave_translator:uav_waitrequest -> lcd_control_slave_translator_avalon_universal_slave_0_agent:m0_waitrequest
	signal lcd_control_slave_translator_avalon_universal_slave_0_agent_m0_burstcount                         : std_logic_vector(2 downto 0);  -- lcd_control_slave_translator_avalon_universal_slave_0_agent:m0_burstcount -> lcd_control_slave_translator:uav_burstcount
	signal lcd_control_slave_translator_avalon_universal_slave_0_agent_m0_writedata                          : std_logic_vector(31 downto 0); -- lcd_control_slave_translator_avalon_universal_slave_0_agent:m0_writedata -> lcd_control_slave_translator:uav_writedata
	signal lcd_control_slave_translator_avalon_universal_slave_0_agent_m0_address                            : std_logic_vector(18 downto 0); -- lcd_control_slave_translator_avalon_universal_slave_0_agent:m0_address -> lcd_control_slave_translator:uav_address
	signal lcd_control_slave_translator_avalon_universal_slave_0_agent_m0_write                              : std_logic;                     -- lcd_control_slave_translator_avalon_universal_slave_0_agent:m0_write -> lcd_control_slave_translator:uav_write
	signal lcd_control_slave_translator_avalon_universal_slave_0_agent_m0_lock                               : std_logic;                     -- lcd_control_slave_translator_avalon_universal_slave_0_agent:m0_lock -> lcd_control_slave_translator:uav_lock
	signal lcd_control_slave_translator_avalon_universal_slave_0_agent_m0_read                               : std_logic;                     -- lcd_control_slave_translator_avalon_universal_slave_0_agent:m0_read -> lcd_control_slave_translator:uav_read
	signal lcd_control_slave_translator_avalon_universal_slave_0_agent_m0_readdata                           : std_logic_vector(31 downto 0); -- lcd_control_slave_translator:uav_readdata -> lcd_control_slave_translator_avalon_universal_slave_0_agent:m0_readdata
	signal lcd_control_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid                      : std_logic;                     -- lcd_control_slave_translator:uav_readdatavalid -> lcd_control_slave_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	signal lcd_control_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess                        : std_logic;                     -- lcd_control_slave_translator_avalon_universal_slave_0_agent:m0_debugaccess -> lcd_control_slave_translator:uav_debugaccess
	signal lcd_control_slave_translator_avalon_universal_slave_0_agent_m0_byteenable                         : std_logic_vector(3 downto 0);  -- lcd_control_slave_translator_avalon_universal_slave_0_agent:m0_byteenable -> lcd_control_slave_translator:uav_byteenable
	signal lcd_control_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket                 : std_logic;                     -- lcd_control_slave_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> lcd_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	signal lcd_control_slave_translator_avalon_universal_slave_0_agent_rf_source_valid                       : std_logic;                     -- lcd_control_slave_translator_avalon_universal_slave_0_agent:rf_source_valid -> lcd_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	signal lcd_control_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket               : std_logic;                     -- lcd_control_slave_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> lcd_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	signal lcd_control_slave_translator_avalon_universal_slave_0_agent_rf_source_data                        : std_logic_vector(76 downto 0); -- lcd_control_slave_translator_avalon_universal_slave_0_agent:rf_source_data -> lcd_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	signal lcd_control_slave_translator_avalon_universal_slave_0_agent_rf_source_ready                       : std_logic;                     -- lcd_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> lcd_control_slave_translator_avalon_universal_slave_0_agent:rf_source_ready
	signal lcd_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket              : std_logic;                     -- lcd_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> lcd_control_slave_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	signal lcd_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid                    : std_logic;                     -- lcd_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> lcd_control_slave_translator_avalon_universal_slave_0_agent:rf_sink_valid
	signal lcd_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket            : std_logic;                     -- lcd_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> lcd_control_slave_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	signal lcd_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data                     : std_logic_vector(76 downto 0); -- lcd_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> lcd_control_slave_translator_avalon_universal_slave_0_agent:rf_sink_data
	signal lcd_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready                    : std_logic;                     -- lcd_control_slave_translator_avalon_universal_slave_0_agent:rf_sink_ready -> lcd_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	signal lcd_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid                  : std_logic;                     -- lcd_control_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> lcd_control_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	signal lcd_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data                   : std_logic_vector(31 downto 0); -- lcd_control_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> lcd_control_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	signal lcd_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready                  : std_logic;                     -- lcd_control_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> lcd_control_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	signal nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_waitrequest             : std_logic;                     -- nios2_qsys_jtag_debug_module_translator:uav_waitrequest -> nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_waitrequest
	signal nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_burstcount              : std_logic_vector(2 downto 0);  -- nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_burstcount -> nios2_qsys_jtag_debug_module_translator:uav_burstcount
	signal nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_writedata               : std_logic_vector(31 downto 0); -- nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_writedata -> nios2_qsys_jtag_debug_module_translator:uav_writedata
	signal nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_address                 : std_logic_vector(18 downto 0); -- nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_address -> nios2_qsys_jtag_debug_module_translator:uav_address
	signal nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_write                   : std_logic;                     -- nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_write -> nios2_qsys_jtag_debug_module_translator:uav_write
	signal nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_lock                    : std_logic;                     -- nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_lock -> nios2_qsys_jtag_debug_module_translator:uav_lock
	signal nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_read                    : std_logic;                     -- nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_read -> nios2_qsys_jtag_debug_module_translator:uav_read
	signal nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_readdata                : std_logic_vector(31 downto 0); -- nios2_qsys_jtag_debug_module_translator:uav_readdata -> nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_readdata
	signal nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_readdatavalid           : std_logic;                     -- nios2_qsys_jtag_debug_module_translator:uav_readdatavalid -> nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	signal nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_debugaccess             : std_logic;                     -- nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_debugaccess -> nios2_qsys_jtag_debug_module_translator:uav_debugaccess
	signal nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_byteenable              : std_logic_vector(3 downto 0);  -- nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_byteenable -> nios2_qsys_jtag_debug_module_translator:uav_byteenable
	signal nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_endofpacket      : std_logic;                     -- nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	signal nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_valid            : std_logic;                     -- nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_source_valid -> nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	signal nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_startofpacket    : std_logic;                     -- nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	signal nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_data             : std_logic_vector(76 downto 0); -- nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_source_data -> nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	signal nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_ready            : std_logic;                     -- nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_source_ready
	signal nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket   : std_logic;                     -- nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	signal nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid         : std_logic;                     -- nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_sink_valid
	signal nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket : std_logic;                     -- nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	signal nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data          : std_logic_vector(76 downto 0); -- nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_sink_data
	signal nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready         : std_logic;                     -- nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_sink_ready -> nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	signal nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid       : std_logic;                     -- nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	signal nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data        : std_logic_vector(31 downto 0); -- nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	signal nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready       : std_logic;                     -- nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	signal nios2_qsys_instruction_master_translator_avalon_universal_master_0_waitrequest                    : std_logic;                     -- nios2_qsys_instruction_master_translator_avalon_universal_master_0_agent:av_waitrequest -> nios2_qsys_instruction_master_translator:uav_waitrequest
	signal nios2_qsys_instruction_master_translator_avalon_universal_master_0_burstcount                     : std_logic_vector(2 downto 0);  -- nios2_qsys_instruction_master_translator:uav_burstcount -> nios2_qsys_instruction_master_translator_avalon_universal_master_0_agent:av_burstcount
	signal nios2_qsys_instruction_master_translator_avalon_universal_master_0_writedata                      : std_logic_vector(31 downto 0); -- nios2_qsys_instruction_master_translator:uav_writedata -> nios2_qsys_instruction_master_translator_avalon_universal_master_0_agent:av_writedata
	signal nios2_qsys_instruction_master_translator_avalon_universal_master_0_address                        : std_logic_vector(18 downto 0); -- nios2_qsys_instruction_master_translator:uav_address -> nios2_qsys_instruction_master_translator_avalon_universal_master_0_agent:av_address
	signal nios2_qsys_instruction_master_translator_avalon_universal_master_0_lock                           : std_logic;                     -- nios2_qsys_instruction_master_translator:uav_lock -> nios2_qsys_instruction_master_translator_avalon_universal_master_0_agent:av_lock
	signal nios2_qsys_instruction_master_translator_avalon_universal_master_0_write                          : std_logic;                     -- nios2_qsys_instruction_master_translator:uav_write -> nios2_qsys_instruction_master_translator_avalon_universal_master_0_agent:av_write
	signal nios2_qsys_instruction_master_translator_avalon_universal_master_0_read                           : std_logic;                     -- nios2_qsys_instruction_master_translator:uav_read -> nios2_qsys_instruction_master_translator_avalon_universal_master_0_agent:av_read
	signal nios2_qsys_instruction_master_translator_avalon_universal_master_0_readdata                       : std_logic_vector(31 downto 0); -- nios2_qsys_instruction_master_translator_avalon_universal_master_0_agent:av_readdata -> nios2_qsys_instruction_master_translator:uav_readdata
	signal nios2_qsys_instruction_master_translator_avalon_universal_master_0_debugaccess                    : std_logic;                     -- nios2_qsys_instruction_master_translator:uav_debugaccess -> nios2_qsys_instruction_master_translator_avalon_universal_master_0_agent:av_debugaccess
	signal nios2_qsys_instruction_master_translator_avalon_universal_master_0_byteenable                     : std_logic_vector(3 downto 0);  -- nios2_qsys_instruction_master_translator:uav_byteenable -> nios2_qsys_instruction_master_translator_avalon_universal_master_0_agent:av_byteenable
	signal nios2_qsys_instruction_master_translator_avalon_universal_master_0_readdatavalid                  : std_logic;                     -- nios2_qsys_instruction_master_translator_avalon_universal_master_0_agent:av_readdatavalid -> nios2_qsys_instruction_master_translator:uav_readdatavalid
	signal pio_sw_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest                                : std_logic;                     -- pio_SW_s1_translator:uav_waitrequest -> pio_SW_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	signal pio_sw_s1_translator_avalon_universal_slave_0_agent_m0_burstcount                                 : std_logic_vector(2 downto 0);  -- pio_SW_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> pio_SW_s1_translator:uav_burstcount
	signal pio_sw_s1_translator_avalon_universal_slave_0_agent_m0_writedata                                  : std_logic_vector(31 downto 0); -- pio_SW_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> pio_SW_s1_translator:uav_writedata
	signal pio_sw_s1_translator_avalon_universal_slave_0_agent_m0_address                                    : std_logic_vector(18 downto 0); -- pio_SW_s1_translator_avalon_universal_slave_0_agent:m0_address -> pio_SW_s1_translator:uav_address
	signal pio_sw_s1_translator_avalon_universal_slave_0_agent_m0_write                                      : std_logic;                     -- pio_SW_s1_translator_avalon_universal_slave_0_agent:m0_write -> pio_SW_s1_translator:uav_write
	signal pio_sw_s1_translator_avalon_universal_slave_0_agent_m0_lock                                       : std_logic;                     -- pio_SW_s1_translator_avalon_universal_slave_0_agent:m0_lock -> pio_SW_s1_translator:uav_lock
	signal pio_sw_s1_translator_avalon_universal_slave_0_agent_m0_read                                       : std_logic;                     -- pio_SW_s1_translator_avalon_universal_slave_0_agent:m0_read -> pio_SW_s1_translator:uav_read
	signal pio_sw_s1_translator_avalon_universal_slave_0_agent_m0_readdata                                   : std_logic_vector(31 downto 0); -- pio_SW_s1_translator:uav_readdata -> pio_SW_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	signal pio_sw_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid                              : std_logic;                     -- pio_SW_s1_translator:uav_readdatavalid -> pio_SW_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	signal pio_sw_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess                                : std_logic;                     -- pio_SW_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> pio_SW_s1_translator:uav_debugaccess
	signal pio_sw_s1_translator_avalon_universal_slave_0_agent_m0_byteenable                                 : std_logic_vector(3 downto 0);  -- pio_SW_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> pio_SW_s1_translator:uav_byteenable
	signal pio_sw_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket                         : std_logic;                     -- pio_SW_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> pio_SW_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	signal pio_sw_s1_translator_avalon_universal_slave_0_agent_rf_source_valid                               : std_logic;                     -- pio_SW_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> pio_SW_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	signal pio_sw_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket                       : std_logic;                     -- pio_SW_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> pio_SW_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	signal pio_sw_s1_translator_avalon_universal_slave_0_agent_rf_source_data                                : std_logic_vector(76 downto 0); -- pio_SW_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> pio_SW_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	signal pio_sw_s1_translator_avalon_universal_slave_0_agent_rf_source_ready                               : std_logic;                     -- pio_SW_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> pio_SW_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	signal pio_sw_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket                      : std_logic;                     -- pio_SW_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> pio_SW_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	signal pio_sw_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid                            : std_logic;                     -- pio_SW_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> pio_SW_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	signal pio_sw_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket                    : std_logic;                     -- pio_SW_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> pio_SW_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	signal pio_sw_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data                             : std_logic_vector(76 downto 0); -- pio_SW_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> pio_SW_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	signal pio_sw_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready                            : std_logic;                     -- pio_SW_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> pio_SW_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	signal pio_sw_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid                          : std_logic;                     -- pio_SW_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> pio_SW_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	signal pio_sw_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data                           : std_logic_vector(31 downto 0); -- pio_SW_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> pio_SW_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	signal pio_sw_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready                          : std_logic;                     -- pio_SW_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> pio_SW_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	signal jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest              : std_logic;                     -- jtag_uart_avalon_jtag_slave_translator:uav_waitrequest -> jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_waitrequest
	signal jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_burstcount               : std_logic_vector(2 downto 0);  -- jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_burstcount -> jtag_uart_avalon_jtag_slave_translator:uav_burstcount
	signal jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_writedata                : std_logic_vector(31 downto 0); -- jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_writedata -> jtag_uart_avalon_jtag_slave_translator:uav_writedata
	signal jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_address                  : std_logic_vector(18 downto 0); -- jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_address -> jtag_uart_avalon_jtag_slave_translator:uav_address
	signal jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_write                    : std_logic;                     -- jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_write -> jtag_uart_avalon_jtag_slave_translator:uav_write
	signal jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_lock                     : std_logic;                     -- jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_lock -> jtag_uart_avalon_jtag_slave_translator:uav_lock
	signal jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_read                     : std_logic;                     -- jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_read -> jtag_uart_avalon_jtag_slave_translator:uav_read
	signal jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_readdata                 : std_logic_vector(31 downto 0); -- jtag_uart_avalon_jtag_slave_translator:uav_readdata -> jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_readdata
	signal jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid            : std_logic;                     -- jtag_uart_avalon_jtag_slave_translator:uav_readdatavalid -> jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	signal jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess              : std_logic;                     -- jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_debugaccess -> jtag_uart_avalon_jtag_slave_translator:uav_debugaccess
	signal jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_byteenable               : std_logic_vector(3 downto 0);  -- jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_byteenable -> jtag_uart_avalon_jtag_slave_translator:uav_byteenable
	signal jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket       : std_logic;                     -- jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	signal jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_valid             : std_logic;                     -- jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_source_valid -> jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	signal jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket     : std_logic;                     -- jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	signal jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_data              : std_logic_vector(76 downto 0); -- jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_source_data -> jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	signal jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_ready             : std_logic;                     -- jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_source_ready
	signal jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket    : std_logic;                     -- jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	signal jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid          : std_logic;                     -- jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_sink_valid
	signal jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket  : std_logic;                     -- jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	signal jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data           : std_logic_vector(76 downto 0); -- jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_sink_data
	signal jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready          : std_logic;                     -- jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_sink_ready -> jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	signal jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid        : std_logic;                     -- jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	signal jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data         : std_logic_vector(31 downto 0); -- jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	signal jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready        : std_logic;                     -- jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	signal pio_button_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest                            : std_logic;                     -- pio_Button_s1_translator:uav_waitrequest -> pio_Button_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	signal pio_button_s1_translator_avalon_universal_slave_0_agent_m0_burstcount                             : std_logic_vector(2 downto 0);  -- pio_Button_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> pio_Button_s1_translator:uav_burstcount
	signal pio_button_s1_translator_avalon_universal_slave_0_agent_m0_writedata                              : std_logic_vector(31 downto 0); -- pio_Button_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> pio_Button_s1_translator:uav_writedata
	signal pio_button_s1_translator_avalon_universal_slave_0_agent_m0_address                                : std_logic_vector(18 downto 0); -- pio_Button_s1_translator_avalon_universal_slave_0_agent:m0_address -> pio_Button_s1_translator:uav_address
	signal pio_button_s1_translator_avalon_universal_slave_0_agent_m0_write                                  : std_logic;                     -- pio_Button_s1_translator_avalon_universal_slave_0_agent:m0_write -> pio_Button_s1_translator:uav_write
	signal pio_button_s1_translator_avalon_universal_slave_0_agent_m0_lock                                   : std_logic;                     -- pio_Button_s1_translator_avalon_universal_slave_0_agent:m0_lock -> pio_Button_s1_translator:uav_lock
	signal pio_button_s1_translator_avalon_universal_slave_0_agent_m0_read                                   : std_logic;                     -- pio_Button_s1_translator_avalon_universal_slave_0_agent:m0_read -> pio_Button_s1_translator:uav_read
	signal pio_button_s1_translator_avalon_universal_slave_0_agent_m0_readdata                               : std_logic_vector(31 downto 0); -- pio_Button_s1_translator:uav_readdata -> pio_Button_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	signal pio_button_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid                          : std_logic;                     -- pio_Button_s1_translator:uav_readdatavalid -> pio_Button_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	signal pio_button_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess                            : std_logic;                     -- pio_Button_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> pio_Button_s1_translator:uav_debugaccess
	signal pio_button_s1_translator_avalon_universal_slave_0_agent_m0_byteenable                             : std_logic_vector(3 downto 0);  -- pio_Button_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> pio_Button_s1_translator:uav_byteenable
	signal pio_button_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket                     : std_logic;                     -- pio_Button_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> pio_Button_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	signal pio_button_s1_translator_avalon_universal_slave_0_agent_rf_source_valid                           : std_logic;                     -- pio_Button_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> pio_Button_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	signal pio_button_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket                   : std_logic;                     -- pio_Button_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> pio_Button_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	signal pio_button_s1_translator_avalon_universal_slave_0_agent_rf_source_data                            : std_logic_vector(76 downto 0); -- pio_Button_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> pio_Button_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	signal pio_button_s1_translator_avalon_universal_slave_0_agent_rf_source_ready                           : std_logic;                     -- pio_Button_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> pio_Button_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	signal pio_button_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket                  : std_logic;                     -- pio_Button_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> pio_Button_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	signal pio_button_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid                        : std_logic;                     -- pio_Button_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> pio_Button_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	signal pio_button_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket                : std_logic;                     -- pio_Button_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> pio_Button_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	signal pio_button_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data                         : std_logic_vector(76 downto 0); -- pio_Button_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> pio_Button_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	signal pio_button_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready                        : std_logic;                     -- pio_Button_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> pio_Button_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	signal pio_button_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid                      : std_logic;                     -- pio_Button_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> pio_Button_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	signal pio_button_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data                       : std_logic_vector(31 downto 0); -- pio_Button_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> pio_Button_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	signal pio_button_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready                      : std_logic;                     -- pio_Button_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> pio_Button_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	signal pio_data_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest                              : std_logic;                     -- pio_Data_s1_translator:uav_waitrequest -> pio_Data_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	signal pio_data_s1_translator_avalon_universal_slave_0_agent_m0_burstcount                               : std_logic_vector(2 downto 0);  -- pio_Data_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> pio_Data_s1_translator:uav_burstcount
	signal pio_data_s1_translator_avalon_universal_slave_0_agent_m0_writedata                                : std_logic_vector(31 downto 0); -- pio_Data_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> pio_Data_s1_translator:uav_writedata
	signal pio_data_s1_translator_avalon_universal_slave_0_agent_m0_address                                  : std_logic_vector(18 downto 0); -- pio_Data_s1_translator_avalon_universal_slave_0_agent:m0_address -> pio_Data_s1_translator:uav_address
	signal pio_data_s1_translator_avalon_universal_slave_0_agent_m0_write                                    : std_logic;                     -- pio_Data_s1_translator_avalon_universal_slave_0_agent:m0_write -> pio_Data_s1_translator:uav_write
	signal pio_data_s1_translator_avalon_universal_slave_0_agent_m0_lock                                     : std_logic;                     -- pio_Data_s1_translator_avalon_universal_slave_0_agent:m0_lock -> pio_Data_s1_translator:uav_lock
	signal pio_data_s1_translator_avalon_universal_slave_0_agent_m0_read                                     : std_logic;                     -- pio_Data_s1_translator_avalon_universal_slave_0_agent:m0_read -> pio_Data_s1_translator:uav_read
	signal pio_data_s1_translator_avalon_universal_slave_0_agent_m0_readdata                                 : std_logic_vector(31 downto 0); -- pio_Data_s1_translator:uav_readdata -> pio_Data_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	signal pio_data_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid                            : std_logic;                     -- pio_Data_s1_translator:uav_readdatavalid -> pio_Data_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	signal pio_data_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess                              : std_logic;                     -- pio_Data_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> pio_Data_s1_translator:uav_debugaccess
	signal pio_data_s1_translator_avalon_universal_slave_0_agent_m0_byteenable                               : std_logic_vector(3 downto 0);  -- pio_Data_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> pio_Data_s1_translator:uav_byteenable
	signal pio_data_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket                       : std_logic;                     -- pio_Data_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> pio_Data_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	signal pio_data_s1_translator_avalon_universal_slave_0_agent_rf_source_valid                             : std_logic;                     -- pio_Data_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> pio_Data_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	signal pio_data_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket                     : std_logic;                     -- pio_Data_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> pio_Data_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	signal pio_data_s1_translator_avalon_universal_slave_0_agent_rf_source_data                              : std_logic_vector(76 downto 0); -- pio_Data_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> pio_Data_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	signal pio_data_s1_translator_avalon_universal_slave_0_agent_rf_source_ready                             : std_logic;                     -- pio_Data_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> pio_Data_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	signal pio_data_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket                    : std_logic;                     -- pio_Data_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> pio_Data_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	signal pio_data_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid                          : std_logic;                     -- pio_Data_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> pio_Data_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	signal pio_data_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket                  : std_logic;                     -- pio_Data_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> pio_Data_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	signal pio_data_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data                           : std_logic_vector(76 downto 0); -- pio_Data_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> pio_Data_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	signal pio_data_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready                          : std_logic;                     -- pio_Data_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> pio_Data_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	signal pio_data_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid                        : std_logic;                     -- pio_Data_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> pio_Data_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	signal pio_data_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data                         : std_logic_vector(31 downto 0); -- pio_Data_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> pio_Data_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	signal pio_data_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready                        : std_logic;                     -- pio_Data_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> pio_Data_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	signal uart_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest                                  : std_logic;                     -- uart_s1_translator:uav_waitrequest -> uart_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	signal uart_s1_translator_avalon_universal_slave_0_agent_m0_burstcount                                   : std_logic_vector(2 downto 0);  -- uart_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> uart_s1_translator:uav_burstcount
	signal uart_s1_translator_avalon_universal_slave_0_agent_m0_writedata                                    : std_logic_vector(31 downto 0); -- uart_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> uart_s1_translator:uav_writedata
	signal uart_s1_translator_avalon_universal_slave_0_agent_m0_address                                      : std_logic_vector(18 downto 0); -- uart_s1_translator_avalon_universal_slave_0_agent:m0_address -> uart_s1_translator:uav_address
	signal uart_s1_translator_avalon_universal_slave_0_agent_m0_write                                        : std_logic;                     -- uart_s1_translator_avalon_universal_slave_0_agent:m0_write -> uart_s1_translator:uav_write
	signal uart_s1_translator_avalon_universal_slave_0_agent_m0_lock                                         : std_logic;                     -- uart_s1_translator_avalon_universal_slave_0_agent:m0_lock -> uart_s1_translator:uav_lock
	signal uart_s1_translator_avalon_universal_slave_0_agent_m0_read                                         : std_logic;                     -- uart_s1_translator_avalon_universal_slave_0_agent:m0_read -> uart_s1_translator:uav_read
	signal uart_s1_translator_avalon_universal_slave_0_agent_m0_readdata                                     : std_logic_vector(31 downto 0); -- uart_s1_translator:uav_readdata -> uart_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	signal uart_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid                                : std_logic;                     -- uart_s1_translator:uav_readdatavalid -> uart_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	signal uart_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess                                  : std_logic;                     -- uart_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> uart_s1_translator:uav_debugaccess
	signal uart_s1_translator_avalon_universal_slave_0_agent_m0_byteenable                                   : std_logic_vector(3 downto 0);  -- uart_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> uart_s1_translator:uav_byteenable
	signal uart_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket                           : std_logic;                     -- uart_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> uart_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	signal uart_s1_translator_avalon_universal_slave_0_agent_rf_source_valid                                 : std_logic;                     -- uart_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> uart_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	signal uart_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket                         : std_logic;                     -- uart_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> uart_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	signal uart_s1_translator_avalon_universal_slave_0_agent_rf_source_data                                  : std_logic_vector(76 downto 0); -- uart_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> uart_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	signal uart_s1_translator_avalon_universal_slave_0_agent_rf_source_ready                                 : std_logic;                     -- uart_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> uart_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	signal uart_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket                        : std_logic;                     -- uart_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> uart_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	signal uart_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid                              : std_logic;                     -- uart_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> uart_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	signal uart_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket                      : std_logic;                     -- uart_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> uart_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	signal uart_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data                               : std_logic_vector(76 downto 0); -- uart_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> uart_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	signal uart_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready                              : std_logic;                     -- uart_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> uart_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	signal uart_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid                            : std_logic;                     -- uart_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> uart_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	signal uart_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data                             : std_logic_vector(31 downto 0); -- uart_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> uart_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	signal uart_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready                            : std_logic;                     -- uart_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> uart_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	signal onchip_memory_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest                         : std_logic;                     -- onchip_memory_s1_translator:uav_waitrequest -> onchip_memory_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	signal onchip_memory_s1_translator_avalon_universal_slave_0_agent_m0_burstcount                          : std_logic_vector(2 downto 0);  -- onchip_memory_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> onchip_memory_s1_translator:uav_burstcount
	signal onchip_memory_s1_translator_avalon_universal_slave_0_agent_m0_writedata                           : std_logic_vector(31 downto 0); -- onchip_memory_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> onchip_memory_s1_translator:uav_writedata
	signal onchip_memory_s1_translator_avalon_universal_slave_0_agent_m0_address                             : std_logic_vector(18 downto 0); -- onchip_memory_s1_translator_avalon_universal_slave_0_agent:m0_address -> onchip_memory_s1_translator:uav_address
	signal onchip_memory_s1_translator_avalon_universal_slave_0_agent_m0_write                               : std_logic;                     -- onchip_memory_s1_translator_avalon_universal_slave_0_agent:m0_write -> onchip_memory_s1_translator:uav_write
	signal onchip_memory_s1_translator_avalon_universal_slave_0_agent_m0_lock                                : std_logic;                     -- onchip_memory_s1_translator_avalon_universal_slave_0_agent:m0_lock -> onchip_memory_s1_translator:uav_lock
	signal onchip_memory_s1_translator_avalon_universal_slave_0_agent_m0_read                                : std_logic;                     -- onchip_memory_s1_translator_avalon_universal_slave_0_agent:m0_read -> onchip_memory_s1_translator:uav_read
	signal onchip_memory_s1_translator_avalon_universal_slave_0_agent_m0_readdata                            : std_logic_vector(31 downto 0); -- onchip_memory_s1_translator:uav_readdata -> onchip_memory_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	signal onchip_memory_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid                       : std_logic;                     -- onchip_memory_s1_translator:uav_readdatavalid -> onchip_memory_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	signal onchip_memory_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess                         : std_logic;                     -- onchip_memory_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> onchip_memory_s1_translator:uav_debugaccess
	signal onchip_memory_s1_translator_avalon_universal_slave_0_agent_m0_byteenable                          : std_logic_vector(3 downto 0);  -- onchip_memory_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> onchip_memory_s1_translator:uav_byteenable
	signal onchip_memory_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket                  : std_logic;                     -- onchip_memory_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> onchip_memory_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	signal onchip_memory_s1_translator_avalon_universal_slave_0_agent_rf_source_valid                        : std_logic;                     -- onchip_memory_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> onchip_memory_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	signal onchip_memory_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket                : std_logic;                     -- onchip_memory_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> onchip_memory_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	signal onchip_memory_s1_translator_avalon_universal_slave_0_agent_rf_source_data                         : std_logic_vector(76 downto 0); -- onchip_memory_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> onchip_memory_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	signal onchip_memory_s1_translator_avalon_universal_slave_0_agent_rf_source_ready                        : std_logic;                     -- onchip_memory_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> onchip_memory_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	signal onchip_memory_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket               : std_logic;                     -- onchip_memory_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> onchip_memory_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	signal onchip_memory_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid                     : std_logic;                     -- onchip_memory_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> onchip_memory_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	signal onchip_memory_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket             : std_logic;                     -- onchip_memory_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> onchip_memory_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	signal onchip_memory_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data                      : std_logic_vector(76 downto 0); -- onchip_memory_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> onchip_memory_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	signal onchip_memory_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready                     : std_logic;                     -- onchip_memory_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> onchip_memory_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	signal onchip_memory_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid                   : std_logic;                     -- onchip_memory_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> onchip_memory_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	signal onchip_memory_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data                    : std_logic_vector(31 downto 0); -- onchip_memory_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> onchip_memory_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	signal onchip_memory_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready                   : std_logic;                     -- onchip_memory_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> onchip_memory_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	signal timer_0_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest                               : std_logic;                     -- timer_0_s1_translator:uav_waitrequest -> timer_0_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	signal timer_0_s1_translator_avalon_universal_slave_0_agent_m0_burstcount                                : std_logic_vector(2 downto 0);  -- timer_0_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> timer_0_s1_translator:uav_burstcount
	signal timer_0_s1_translator_avalon_universal_slave_0_agent_m0_writedata                                 : std_logic_vector(31 downto 0); -- timer_0_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> timer_0_s1_translator:uav_writedata
	signal timer_0_s1_translator_avalon_universal_slave_0_agent_m0_address                                   : std_logic_vector(18 downto 0); -- timer_0_s1_translator_avalon_universal_slave_0_agent:m0_address -> timer_0_s1_translator:uav_address
	signal timer_0_s1_translator_avalon_universal_slave_0_agent_m0_write                                     : std_logic;                     -- timer_0_s1_translator_avalon_universal_slave_0_agent:m0_write -> timer_0_s1_translator:uav_write
	signal timer_0_s1_translator_avalon_universal_slave_0_agent_m0_lock                                      : std_logic;                     -- timer_0_s1_translator_avalon_universal_slave_0_agent:m0_lock -> timer_0_s1_translator:uav_lock
	signal timer_0_s1_translator_avalon_universal_slave_0_agent_m0_read                                      : std_logic;                     -- timer_0_s1_translator_avalon_universal_slave_0_agent:m0_read -> timer_0_s1_translator:uav_read
	signal timer_0_s1_translator_avalon_universal_slave_0_agent_m0_readdata                                  : std_logic_vector(31 downto 0); -- timer_0_s1_translator:uav_readdata -> timer_0_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	signal timer_0_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid                             : std_logic;                     -- timer_0_s1_translator:uav_readdatavalid -> timer_0_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	signal timer_0_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess                               : std_logic;                     -- timer_0_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> timer_0_s1_translator:uav_debugaccess
	signal timer_0_s1_translator_avalon_universal_slave_0_agent_m0_byteenable                                : std_logic_vector(3 downto 0);  -- timer_0_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> timer_0_s1_translator:uav_byteenable
	signal timer_0_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket                        : std_logic;                     -- timer_0_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> timer_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	signal timer_0_s1_translator_avalon_universal_slave_0_agent_rf_source_valid                              : std_logic;                     -- timer_0_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> timer_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	signal timer_0_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket                      : std_logic;                     -- timer_0_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> timer_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	signal timer_0_s1_translator_avalon_universal_slave_0_agent_rf_source_data                               : std_logic_vector(76 downto 0); -- timer_0_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> timer_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	signal timer_0_s1_translator_avalon_universal_slave_0_agent_rf_source_ready                              : std_logic;                     -- timer_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> timer_0_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	signal timer_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket                     : std_logic;                     -- timer_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> timer_0_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	signal timer_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid                           : std_logic;                     -- timer_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> timer_0_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	signal timer_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket                   : std_logic;                     -- timer_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> timer_0_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	signal timer_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data                            : std_logic_vector(76 downto 0); -- timer_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> timer_0_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	signal timer_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready                           : std_logic;                     -- timer_0_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> timer_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	signal timer_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid                         : std_logic;                     -- timer_0_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> timer_0_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	signal timer_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data                          : std_logic_vector(31 downto 0); -- timer_0_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> timer_0_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	signal timer_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready                         : std_logic;                     -- timer_0_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> timer_0_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	signal pio_rdydata_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest                           : std_logic;                     -- pio_RdyData_s1_translator:uav_waitrequest -> pio_RdyData_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	signal pio_rdydata_s1_translator_avalon_universal_slave_0_agent_m0_burstcount                            : std_logic_vector(2 downto 0);  -- pio_RdyData_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> pio_RdyData_s1_translator:uav_burstcount
	signal pio_rdydata_s1_translator_avalon_universal_slave_0_agent_m0_writedata                             : std_logic_vector(31 downto 0); -- pio_RdyData_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> pio_RdyData_s1_translator:uav_writedata
	signal pio_rdydata_s1_translator_avalon_universal_slave_0_agent_m0_address                               : std_logic_vector(18 downto 0); -- pio_RdyData_s1_translator_avalon_universal_slave_0_agent:m0_address -> pio_RdyData_s1_translator:uav_address
	signal pio_rdydata_s1_translator_avalon_universal_slave_0_agent_m0_write                                 : std_logic;                     -- pio_RdyData_s1_translator_avalon_universal_slave_0_agent:m0_write -> pio_RdyData_s1_translator:uav_write
	signal pio_rdydata_s1_translator_avalon_universal_slave_0_agent_m0_lock                                  : std_logic;                     -- pio_RdyData_s1_translator_avalon_universal_slave_0_agent:m0_lock -> pio_RdyData_s1_translator:uav_lock
	signal pio_rdydata_s1_translator_avalon_universal_slave_0_agent_m0_read                                  : std_logic;                     -- pio_RdyData_s1_translator_avalon_universal_slave_0_agent:m0_read -> pio_RdyData_s1_translator:uav_read
	signal pio_rdydata_s1_translator_avalon_universal_slave_0_agent_m0_readdata                              : std_logic_vector(31 downto 0); -- pio_RdyData_s1_translator:uav_readdata -> pio_RdyData_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	signal pio_rdydata_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid                         : std_logic;                     -- pio_RdyData_s1_translator:uav_readdatavalid -> pio_RdyData_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	signal pio_rdydata_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess                           : std_logic;                     -- pio_RdyData_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> pio_RdyData_s1_translator:uav_debugaccess
	signal pio_rdydata_s1_translator_avalon_universal_slave_0_agent_m0_byteenable                            : std_logic_vector(3 downto 0);  -- pio_RdyData_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> pio_RdyData_s1_translator:uav_byteenable
	signal pio_rdydata_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket                    : std_logic;                     -- pio_RdyData_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> pio_RdyData_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	signal pio_rdydata_s1_translator_avalon_universal_slave_0_agent_rf_source_valid                          : std_logic;                     -- pio_RdyData_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> pio_RdyData_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	signal pio_rdydata_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket                  : std_logic;                     -- pio_RdyData_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> pio_RdyData_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	signal pio_rdydata_s1_translator_avalon_universal_slave_0_agent_rf_source_data                           : std_logic_vector(76 downto 0); -- pio_RdyData_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> pio_RdyData_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	signal pio_rdydata_s1_translator_avalon_universal_slave_0_agent_rf_source_ready                          : std_logic;                     -- pio_RdyData_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> pio_RdyData_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	signal pio_rdydata_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket                 : std_logic;                     -- pio_RdyData_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> pio_RdyData_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	signal pio_rdydata_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid                       : std_logic;                     -- pio_RdyData_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> pio_RdyData_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	signal pio_rdydata_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket               : std_logic;                     -- pio_RdyData_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> pio_RdyData_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	signal pio_rdydata_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data                        : std_logic_vector(76 downto 0); -- pio_RdyData_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> pio_RdyData_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	signal pio_rdydata_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready                       : std_logic;                     -- pio_RdyData_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> pio_RdyData_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	signal pio_rdydata_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid                     : std_logic;                     -- pio_RdyData_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> pio_RdyData_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	signal pio_rdydata_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data                      : std_logic_vector(31 downto 0); -- pio_RdyData_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> pio_RdyData_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	signal pio_rdydata_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready                     : std_logic;                     -- pio_RdyData_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> pio_RdyData_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	signal nios2_qsys_instruction_master_translator_avalon_universal_master_0_agent_cp_endofpacket           : std_logic;                     -- nios2_qsys_instruction_master_translator_avalon_universal_master_0_agent:cp_endofpacket -> addr_router:sink_endofpacket
	signal nios2_qsys_instruction_master_translator_avalon_universal_master_0_agent_cp_valid                 : std_logic;                     -- nios2_qsys_instruction_master_translator_avalon_universal_master_0_agent:cp_valid -> addr_router:sink_valid
	signal nios2_qsys_instruction_master_translator_avalon_universal_master_0_agent_cp_startofpacket         : std_logic;                     -- nios2_qsys_instruction_master_translator_avalon_universal_master_0_agent:cp_startofpacket -> addr_router:sink_startofpacket
	signal nios2_qsys_instruction_master_translator_avalon_universal_master_0_agent_cp_data                  : std_logic_vector(75 downto 0); -- nios2_qsys_instruction_master_translator_avalon_universal_master_0_agent:cp_data -> addr_router:sink_data
	signal nios2_qsys_instruction_master_translator_avalon_universal_master_0_agent_cp_ready                 : std_logic;                     -- addr_router:sink_ready -> nios2_qsys_instruction_master_translator_avalon_universal_master_0_agent:cp_ready
	signal nios2_qsys_data_master_translator_avalon_universal_master_0_agent_cp_endofpacket                  : std_logic;                     -- nios2_qsys_data_master_translator_avalon_universal_master_0_agent:cp_endofpacket -> addr_router_001:sink_endofpacket
	signal nios2_qsys_data_master_translator_avalon_universal_master_0_agent_cp_valid                        : std_logic;                     -- nios2_qsys_data_master_translator_avalon_universal_master_0_agent:cp_valid -> addr_router_001:sink_valid
	signal nios2_qsys_data_master_translator_avalon_universal_master_0_agent_cp_startofpacket                : std_logic;                     -- nios2_qsys_data_master_translator_avalon_universal_master_0_agent:cp_startofpacket -> addr_router_001:sink_startofpacket
	signal nios2_qsys_data_master_translator_avalon_universal_master_0_agent_cp_data                         : std_logic_vector(75 downto 0); -- nios2_qsys_data_master_translator_avalon_universal_master_0_agent:cp_data -> addr_router_001:sink_data
	signal nios2_qsys_data_master_translator_avalon_universal_master_0_agent_cp_ready                        : std_logic;                     -- addr_router_001:sink_ready -> nios2_qsys_data_master_translator_avalon_universal_master_0_agent:cp_ready
	signal nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_endofpacket             : std_logic;                     -- nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router:sink_endofpacket
	signal nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_valid                   : std_logic;                     -- nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent:rp_valid -> id_router:sink_valid
	signal nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_startofpacket           : std_logic;                     -- nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router:sink_startofpacket
	signal nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_data                    : std_logic_vector(75 downto 0); -- nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent:rp_data -> id_router:sink_data
	signal nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_ready                   : std_logic;                     -- id_router:sink_ready -> nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent:rp_ready
	signal onchip_memory_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket                         : std_logic;                     -- onchip_memory_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_001:sink_endofpacket
	signal onchip_memory_s1_translator_avalon_universal_slave_0_agent_rp_valid                               : std_logic;                     -- onchip_memory_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_001:sink_valid
	signal onchip_memory_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket                       : std_logic;                     -- onchip_memory_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_001:sink_startofpacket
	signal onchip_memory_s1_translator_avalon_universal_slave_0_agent_rp_data                                : std_logic_vector(75 downto 0); -- onchip_memory_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_001:sink_data
	signal onchip_memory_s1_translator_avalon_universal_slave_0_agent_rp_ready                               : std_logic;                     -- id_router_001:sink_ready -> onchip_memory_s1_translator_avalon_universal_slave_0_agent:rp_ready
	signal jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket              : std_logic;                     -- jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_002:sink_endofpacket
	signal jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_valid                    : std_logic;                     -- jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_002:sink_valid
	signal jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket            : std_logic;                     -- jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_002:sink_startofpacket
	signal jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_data                     : std_logic_vector(75 downto 0); -- jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rp_data -> id_router_002:sink_data
	signal jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_ready                    : std_logic;                     -- id_router_002:sink_ready -> jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rp_ready
	signal sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket                 : std_logic;                     -- sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_003:sink_endofpacket
	signal sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent_rp_valid                       : std_logic;                     -- sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_003:sink_valid
	signal sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket               : std_logic;                     -- sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_003:sink_startofpacket
	signal sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent_rp_data                        : std_logic_vector(75 downto 0); -- sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent:rp_data -> id_router_003:sink_data
	signal sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent_rp_ready                       : std_logic;                     -- id_router_003:sink_ready -> sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent:rp_ready
	signal pio_ledg_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket                              : std_logic;                     -- pio_LEDG_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_004:sink_endofpacket
	signal pio_ledg_s1_translator_avalon_universal_slave_0_agent_rp_valid                                    : std_logic;                     -- pio_LEDG_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_004:sink_valid
	signal pio_ledg_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket                            : std_logic;                     -- pio_LEDG_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_004:sink_startofpacket
	signal pio_ledg_s1_translator_avalon_universal_slave_0_agent_rp_data                                     : std_logic_vector(75 downto 0); -- pio_LEDG_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_004:sink_data
	signal pio_ledg_s1_translator_avalon_universal_slave_0_agent_rp_ready                                    : std_logic;                     -- id_router_004:sink_ready -> pio_LEDG_s1_translator_avalon_universal_slave_0_agent:rp_ready
	signal pio_ledr_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket                              : std_logic;                     -- pio_LEDR_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_005:sink_endofpacket
	signal pio_ledr_s1_translator_avalon_universal_slave_0_agent_rp_valid                                    : std_logic;                     -- pio_LEDR_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_005:sink_valid
	signal pio_ledr_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket                            : std_logic;                     -- pio_LEDR_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_005:sink_startofpacket
	signal pio_ledr_s1_translator_avalon_universal_slave_0_agent_rp_data                                     : std_logic_vector(75 downto 0); -- pio_LEDR_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_005:sink_data
	signal pio_ledr_s1_translator_avalon_universal_slave_0_agent_rp_ready                                    : std_logic;                     -- id_router_005:sink_ready -> pio_LEDR_s1_translator_avalon_universal_slave_0_agent:rp_ready
	signal pio_sw_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket                                : std_logic;                     -- pio_SW_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_006:sink_endofpacket
	signal pio_sw_s1_translator_avalon_universal_slave_0_agent_rp_valid                                      : std_logic;                     -- pio_SW_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_006:sink_valid
	signal pio_sw_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket                              : std_logic;                     -- pio_SW_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_006:sink_startofpacket
	signal pio_sw_s1_translator_avalon_universal_slave_0_agent_rp_data                                       : std_logic_vector(75 downto 0); -- pio_SW_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_006:sink_data
	signal pio_sw_s1_translator_avalon_universal_slave_0_agent_rp_ready                                      : std_logic;                     -- id_router_006:sink_ready -> pio_SW_s1_translator_avalon_universal_slave_0_agent:rp_ready
	signal pio_button_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket                            : std_logic;                     -- pio_Button_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_007:sink_endofpacket
	signal pio_button_s1_translator_avalon_universal_slave_0_agent_rp_valid                                  : std_logic;                     -- pio_Button_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_007:sink_valid
	signal pio_button_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket                          : std_logic;                     -- pio_Button_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_007:sink_startofpacket
	signal pio_button_s1_translator_avalon_universal_slave_0_agent_rp_data                                   : std_logic_vector(75 downto 0); -- pio_Button_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_007:sink_data
	signal pio_button_s1_translator_avalon_universal_slave_0_agent_rp_ready                                  : std_logic;                     -- id_router_007:sink_ready -> pio_Button_s1_translator_avalon_universal_slave_0_agent:rp_ready
	signal lcd_control_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket                        : std_logic;                     -- lcd_control_slave_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_008:sink_endofpacket
	signal lcd_control_slave_translator_avalon_universal_slave_0_agent_rp_valid                              : std_logic;                     -- lcd_control_slave_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_008:sink_valid
	signal lcd_control_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket                      : std_logic;                     -- lcd_control_slave_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_008:sink_startofpacket
	signal lcd_control_slave_translator_avalon_universal_slave_0_agent_rp_data                               : std_logic_vector(75 downto 0); -- lcd_control_slave_translator_avalon_universal_slave_0_agent:rp_data -> id_router_008:sink_data
	signal lcd_control_slave_translator_avalon_universal_slave_0_agent_rp_ready                              : std_logic;                     -- id_router_008:sink_ready -> lcd_control_slave_translator_avalon_universal_slave_0_agent:rp_ready
	signal uart_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket                                  : std_logic;                     -- uart_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_009:sink_endofpacket
	signal uart_s1_translator_avalon_universal_slave_0_agent_rp_valid                                        : std_logic;                     -- uart_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_009:sink_valid
	signal uart_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket                                : std_logic;                     -- uart_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_009:sink_startofpacket
	signal uart_s1_translator_avalon_universal_slave_0_agent_rp_data                                         : std_logic_vector(75 downto 0); -- uart_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_009:sink_data
	signal uart_s1_translator_avalon_universal_slave_0_agent_rp_ready                                        : std_logic;                     -- id_router_009:sink_ready -> uart_s1_translator_avalon_universal_slave_0_agent:rp_ready
	signal timer_0_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket                               : std_logic;                     -- timer_0_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_010:sink_endofpacket
	signal timer_0_s1_translator_avalon_universal_slave_0_agent_rp_valid                                     : std_logic;                     -- timer_0_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_010:sink_valid
	signal timer_0_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket                             : std_logic;                     -- timer_0_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_010:sink_startofpacket
	signal timer_0_s1_translator_avalon_universal_slave_0_agent_rp_data                                      : std_logic_vector(75 downto 0); -- timer_0_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_010:sink_data
	signal timer_0_s1_translator_avalon_universal_slave_0_agent_rp_ready                                     : std_logic;                     -- id_router_010:sink_ready -> timer_0_s1_translator_avalon_universal_slave_0_agent:rp_ready
	signal pio_data_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket                              : std_logic;                     -- pio_Data_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_011:sink_endofpacket
	signal pio_data_s1_translator_avalon_universal_slave_0_agent_rp_valid                                    : std_logic;                     -- pio_Data_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_011:sink_valid
	signal pio_data_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket                            : std_logic;                     -- pio_Data_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_011:sink_startofpacket
	signal pio_data_s1_translator_avalon_universal_slave_0_agent_rp_data                                     : std_logic_vector(75 downto 0); -- pio_Data_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_011:sink_data
	signal pio_data_s1_translator_avalon_universal_slave_0_agent_rp_ready                                    : std_logic;                     -- id_router_011:sink_ready -> pio_Data_s1_translator_avalon_universal_slave_0_agent:rp_ready
	signal pio_rdydata_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket                           : std_logic;                     -- pio_RdyData_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_012:sink_endofpacket
	signal pio_rdydata_s1_translator_avalon_universal_slave_0_agent_rp_valid                                 : std_logic;                     -- pio_RdyData_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_012:sink_valid
	signal pio_rdydata_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket                         : std_logic;                     -- pio_RdyData_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_012:sink_startofpacket
	signal pio_rdydata_s1_translator_avalon_universal_slave_0_agent_rp_data                                  : std_logic_vector(75 downto 0); -- pio_RdyData_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_012:sink_data
	signal pio_rdydata_s1_translator_avalon_universal_slave_0_agent_rp_ready                                 : std_logic;                     -- id_router_012:sink_ready -> pio_RdyData_s1_translator_avalon_universal_slave_0_agent:rp_ready
	signal pio_dataread_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket                          : std_logic;                     -- pio_DataRead_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_013:sink_endofpacket
	signal pio_dataread_s1_translator_avalon_universal_slave_0_agent_rp_valid                                : std_logic;                     -- pio_DataRead_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_013:sink_valid
	signal pio_dataread_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket                        : std_logic;                     -- pio_DataRead_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_013:sink_startofpacket
	signal pio_dataread_s1_translator_avalon_universal_slave_0_agent_rp_data                                 : std_logic_vector(75 downto 0); -- pio_DataRead_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_013:sink_data
	signal pio_dataread_s1_translator_avalon_universal_slave_0_agent_rp_ready                                : std_logic;                     -- id_router_013:sink_ready -> pio_DataRead_s1_translator_avalon_universal_slave_0_agent:rp_ready
	signal addr_router_src_endofpacket                                                                       : std_logic;                     -- addr_router:src_endofpacket -> limiter:cmd_sink_endofpacket
	signal addr_router_src_valid                                                                             : std_logic;                     -- addr_router:src_valid -> limiter:cmd_sink_valid
	signal addr_router_src_startofpacket                                                                     : std_logic;                     -- addr_router:src_startofpacket -> limiter:cmd_sink_startofpacket
	signal addr_router_src_data                                                                              : std_logic_vector(75 downto 0); -- addr_router:src_data -> limiter:cmd_sink_data
	signal addr_router_src_channel                                                                           : std_logic_vector(13 downto 0); -- addr_router:src_channel -> limiter:cmd_sink_channel
	signal addr_router_src_ready                                                                             : std_logic;                     -- limiter:cmd_sink_ready -> addr_router:src_ready
	signal limiter_rsp_src_endofpacket                                                                       : std_logic;                     -- limiter:rsp_src_endofpacket -> nios2_qsys_instruction_master_translator_avalon_universal_master_0_agent:rp_endofpacket
	signal limiter_rsp_src_valid                                                                             : std_logic;                     -- limiter:rsp_src_valid -> nios2_qsys_instruction_master_translator_avalon_universal_master_0_agent:rp_valid
	signal limiter_rsp_src_startofpacket                                                                     : std_logic;                     -- limiter:rsp_src_startofpacket -> nios2_qsys_instruction_master_translator_avalon_universal_master_0_agent:rp_startofpacket
	signal limiter_rsp_src_data                                                                              : std_logic_vector(75 downto 0); -- limiter:rsp_src_data -> nios2_qsys_instruction_master_translator_avalon_universal_master_0_agent:rp_data
	signal limiter_rsp_src_channel                                                                           : std_logic_vector(13 downto 0); -- limiter:rsp_src_channel -> nios2_qsys_instruction_master_translator_avalon_universal_master_0_agent:rp_channel
	signal limiter_rsp_src_ready                                                                             : std_logic;                     -- nios2_qsys_instruction_master_translator_avalon_universal_master_0_agent:rp_ready -> limiter:rsp_src_ready
	signal addr_router_001_src_endofpacket                                                                   : std_logic;                     -- addr_router_001:src_endofpacket -> limiter_001:cmd_sink_endofpacket
	signal addr_router_001_src_valid                                                                         : std_logic;                     -- addr_router_001:src_valid -> limiter_001:cmd_sink_valid
	signal addr_router_001_src_startofpacket                                                                 : std_logic;                     -- addr_router_001:src_startofpacket -> limiter_001:cmd_sink_startofpacket
	signal addr_router_001_src_data                                                                          : std_logic_vector(75 downto 0); -- addr_router_001:src_data -> limiter_001:cmd_sink_data
	signal addr_router_001_src_channel                                                                       : std_logic_vector(13 downto 0); -- addr_router_001:src_channel -> limiter_001:cmd_sink_channel
	signal addr_router_001_src_ready                                                                         : std_logic;                     -- limiter_001:cmd_sink_ready -> addr_router_001:src_ready
	signal limiter_001_rsp_src_endofpacket                                                                   : std_logic;                     -- limiter_001:rsp_src_endofpacket -> nios2_qsys_data_master_translator_avalon_universal_master_0_agent:rp_endofpacket
	signal limiter_001_rsp_src_valid                                                                         : std_logic;                     -- limiter_001:rsp_src_valid -> nios2_qsys_data_master_translator_avalon_universal_master_0_agent:rp_valid
	signal limiter_001_rsp_src_startofpacket                                                                 : std_logic;                     -- limiter_001:rsp_src_startofpacket -> nios2_qsys_data_master_translator_avalon_universal_master_0_agent:rp_startofpacket
	signal limiter_001_rsp_src_data                                                                          : std_logic_vector(75 downto 0); -- limiter_001:rsp_src_data -> nios2_qsys_data_master_translator_avalon_universal_master_0_agent:rp_data
	signal limiter_001_rsp_src_channel                                                                       : std_logic_vector(13 downto 0); -- limiter_001:rsp_src_channel -> nios2_qsys_data_master_translator_avalon_universal_master_0_agent:rp_channel
	signal limiter_001_rsp_src_ready                                                                         : std_logic;                     -- nios2_qsys_data_master_translator_avalon_universal_master_0_agent:rp_ready -> limiter_001:rsp_src_ready
	signal rst_controller_reset_out_reset                                                                    : std_logic;                     -- rst_controller:reset_out -> [addr_router:reset, addr_router_001:reset, cmd_xbar_demux:reset, cmd_xbar_demux_001:reset, cmd_xbar_mux:reset, cmd_xbar_mux_001:reset, id_router:reset, id_router_001:reset, id_router_002:reset, id_router_003:reset, id_router_004:reset, id_router_005:reset, id_router_006:reset, id_router_007:reset, id_router_008:reset, id_router_009:reset, id_router_010:reset, id_router_011:reset, id_router_012:reset, id_router_013:reset, irq_mapper:reset, jtag_uart_avalon_jtag_slave_translator:reset, jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:reset, jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, lcd_control_slave_translator:reset, lcd_control_slave_translator_avalon_universal_slave_0_agent:reset, lcd_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, limiter:reset, limiter_001:reset, nios2_qsys_data_master_translator:reset, nios2_qsys_data_master_translator_avalon_universal_master_0_agent:reset, nios2_qsys_instruction_master_translator:reset, nios2_qsys_instruction_master_translator_avalon_universal_master_0_agent:reset, nios2_qsys_jtag_debug_module_translator:reset, nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent:reset, nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, onchip_memory:reset, onchip_memory_s1_translator:reset, onchip_memory_s1_translator_avalon_universal_slave_0_agent:reset, onchip_memory_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, pio_Button_s1_translator:reset, pio_Button_s1_translator_avalon_universal_slave_0_agent:reset, pio_Button_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, pio_DataRead_s1_translator:reset, pio_DataRead_s1_translator_avalon_universal_slave_0_agent:reset, pio_DataRead_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, pio_Data_s1_translator:reset, pio_Data_s1_translator_avalon_universal_slave_0_agent:reset, pio_Data_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, pio_LEDG_s1_translator:reset, pio_LEDG_s1_translator_avalon_universal_slave_0_agent:reset, pio_LEDG_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, pio_LEDR_s1_translator:reset, pio_LEDR_s1_translator_avalon_universal_slave_0_agent:reset, pio_LEDR_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, pio_RdyData_s1_translator:reset, pio_RdyData_s1_translator_avalon_universal_slave_0_agent:reset, pio_RdyData_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, pio_SW_s1_translator:reset, pio_SW_s1_translator_avalon_universal_slave_0_agent:reset, pio_SW_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, rsp_xbar_demux:reset, rsp_xbar_demux_001:reset, rsp_xbar_demux_002:reset, rsp_xbar_demux_003:reset, rsp_xbar_demux_004:reset, rsp_xbar_demux_005:reset, rsp_xbar_demux_006:reset, rsp_xbar_demux_007:reset, rsp_xbar_demux_008:reset, rsp_xbar_demux_009:reset, rsp_xbar_demux_010:reset, rsp_xbar_demux_011:reset, rsp_xbar_demux_012:reset, rsp_xbar_demux_013:reset, rsp_xbar_mux:reset, rsp_xbar_mux_001:reset, rst_controller_reset_out_reset:in, sysid_qsys_control_slave_translator:reset, sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent:reset, sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, timer_0_s1_translator:reset, timer_0_s1_translator_avalon_universal_slave_0_agent:reset, timer_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, uart_s1_translator:reset, uart_s1_translator_avalon_universal_slave_0_agent:reset, uart_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset]
	signal cmd_xbar_demux_src0_endofpacket                                                                   : std_logic;                     -- cmd_xbar_demux:src0_endofpacket -> cmd_xbar_mux:sink0_endofpacket
	signal cmd_xbar_demux_src0_valid                                                                         : std_logic;                     -- cmd_xbar_demux:src0_valid -> cmd_xbar_mux:sink0_valid
	signal cmd_xbar_demux_src0_startofpacket                                                                 : std_logic;                     -- cmd_xbar_demux:src0_startofpacket -> cmd_xbar_mux:sink0_startofpacket
	signal cmd_xbar_demux_src0_data                                                                          : std_logic_vector(75 downto 0); -- cmd_xbar_demux:src0_data -> cmd_xbar_mux:sink0_data
	signal cmd_xbar_demux_src0_channel                                                                       : std_logic_vector(13 downto 0); -- cmd_xbar_demux:src0_channel -> cmd_xbar_mux:sink0_channel
	signal cmd_xbar_demux_src0_ready                                                                         : std_logic;                     -- cmd_xbar_mux:sink0_ready -> cmd_xbar_demux:src0_ready
	signal cmd_xbar_demux_src1_endofpacket                                                                   : std_logic;                     -- cmd_xbar_demux:src1_endofpacket -> cmd_xbar_mux_001:sink0_endofpacket
	signal cmd_xbar_demux_src1_valid                                                                         : std_logic;                     -- cmd_xbar_demux:src1_valid -> cmd_xbar_mux_001:sink0_valid
	signal cmd_xbar_demux_src1_startofpacket                                                                 : std_logic;                     -- cmd_xbar_demux:src1_startofpacket -> cmd_xbar_mux_001:sink0_startofpacket
	signal cmd_xbar_demux_src1_data                                                                          : std_logic_vector(75 downto 0); -- cmd_xbar_demux:src1_data -> cmd_xbar_mux_001:sink0_data
	signal cmd_xbar_demux_src1_channel                                                                       : std_logic_vector(13 downto 0); -- cmd_xbar_demux:src1_channel -> cmd_xbar_mux_001:sink0_channel
	signal cmd_xbar_demux_src1_ready                                                                         : std_logic;                     -- cmd_xbar_mux_001:sink0_ready -> cmd_xbar_demux:src1_ready
	signal cmd_xbar_demux_001_src0_endofpacket                                                               : std_logic;                     -- cmd_xbar_demux_001:src0_endofpacket -> cmd_xbar_mux:sink1_endofpacket
	signal cmd_xbar_demux_001_src0_valid                                                                     : std_logic;                     -- cmd_xbar_demux_001:src0_valid -> cmd_xbar_mux:sink1_valid
	signal cmd_xbar_demux_001_src0_startofpacket                                                             : std_logic;                     -- cmd_xbar_demux_001:src0_startofpacket -> cmd_xbar_mux:sink1_startofpacket
	signal cmd_xbar_demux_001_src0_data                                                                      : std_logic_vector(75 downto 0); -- cmd_xbar_demux_001:src0_data -> cmd_xbar_mux:sink1_data
	signal cmd_xbar_demux_001_src0_channel                                                                   : std_logic_vector(13 downto 0); -- cmd_xbar_demux_001:src0_channel -> cmd_xbar_mux:sink1_channel
	signal cmd_xbar_demux_001_src0_ready                                                                     : std_logic;                     -- cmd_xbar_mux:sink1_ready -> cmd_xbar_demux_001:src0_ready
	signal cmd_xbar_demux_001_src1_endofpacket                                                               : std_logic;                     -- cmd_xbar_demux_001:src1_endofpacket -> cmd_xbar_mux_001:sink1_endofpacket
	signal cmd_xbar_demux_001_src1_valid                                                                     : std_logic;                     -- cmd_xbar_demux_001:src1_valid -> cmd_xbar_mux_001:sink1_valid
	signal cmd_xbar_demux_001_src1_startofpacket                                                             : std_logic;                     -- cmd_xbar_demux_001:src1_startofpacket -> cmd_xbar_mux_001:sink1_startofpacket
	signal cmd_xbar_demux_001_src1_data                                                                      : std_logic_vector(75 downto 0); -- cmd_xbar_demux_001:src1_data -> cmd_xbar_mux_001:sink1_data
	signal cmd_xbar_demux_001_src1_channel                                                                   : std_logic_vector(13 downto 0); -- cmd_xbar_demux_001:src1_channel -> cmd_xbar_mux_001:sink1_channel
	signal cmd_xbar_demux_001_src1_ready                                                                     : std_logic;                     -- cmd_xbar_mux_001:sink1_ready -> cmd_xbar_demux_001:src1_ready
	signal cmd_xbar_demux_001_src2_endofpacket                                                               : std_logic;                     -- cmd_xbar_demux_001:src2_endofpacket -> jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:cp_endofpacket
	signal cmd_xbar_demux_001_src2_valid                                                                     : std_logic;                     -- cmd_xbar_demux_001:src2_valid -> jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:cp_valid
	signal cmd_xbar_demux_001_src2_startofpacket                                                             : std_logic;                     -- cmd_xbar_demux_001:src2_startofpacket -> jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:cp_startofpacket
	signal cmd_xbar_demux_001_src2_data                                                                      : std_logic_vector(75 downto 0); -- cmd_xbar_demux_001:src2_data -> jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:cp_data
	signal cmd_xbar_demux_001_src2_channel                                                                   : std_logic_vector(13 downto 0); -- cmd_xbar_demux_001:src2_channel -> jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:cp_channel
	signal cmd_xbar_demux_001_src3_endofpacket                                                               : std_logic;                     -- cmd_xbar_demux_001:src3_endofpacket -> sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent:cp_endofpacket
	signal cmd_xbar_demux_001_src3_valid                                                                     : std_logic;                     -- cmd_xbar_demux_001:src3_valid -> sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent:cp_valid
	signal cmd_xbar_demux_001_src3_startofpacket                                                             : std_logic;                     -- cmd_xbar_demux_001:src3_startofpacket -> sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent:cp_startofpacket
	signal cmd_xbar_demux_001_src3_data                                                                      : std_logic_vector(75 downto 0); -- cmd_xbar_demux_001:src3_data -> sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent:cp_data
	signal cmd_xbar_demux_001_src3_channel                                                                   : std_logic_vector(13 downto 0); -- cmd_xbar_demux_001:src3_channel -> sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent:cp_channel
	signal cmd_xbar_demux_001_src4_endofpacket                                                               : std_logic;                     -- cmd_xbar_demux_001:src4_endofpacket -> pio_LEDG_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	signal cmd_xbar_demux_001_src4_valid                                                                     : std_logic;                     -- cmd_xbar_demux_001:src4_valid -> pio_LEDG_s1_translator_avalon_universal_slave_0_agent:cp_valid
	signal cmd_xbar_demux_001_src4_startofpacket                                                             : std_logic;                     -- cmd_xbar_demux_001:src4_startofpacket -> pio_LEDG_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	signal cmd_xbar_demux_001_src4_data                                                                      : std_logic_vector(75 downto 0); -- cmd_xbar_demux_001:src4_data -> pio_LEDG_s1_translator_avalon_universal_slave_0_agent:cp_data
	signal cmd_xbar_demux_001_src4_channel                                                                   : std_logic_vector(13 downto 0); -- cmd_xbar_demux_001:src4_channel -> pio_LEDG_s1_translator_avalon_universal_slave_0_agent:cp_channel
	signal cmd_xbar_demux_001_src5_endofpacket                                                               : std_logic;                     -- cmd_xbar_demux_001:src5_endofpacket -> pio_LEDR_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	signal cmd_xbar_demux_001_src5_valid                                                                     : std_logic;                     -- cmd_xbar_demux_001:src5_valid -> pio_LEDR_s1_translator_avalon_universal_slave_0_agent:cp_valid
	signal cmd_xbar_demux_001_src5_startofpacket                                                             : std_logic;                     -- cmd_xbar_demux_001:src5_startofpacket -> pio_LEDR_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	signal cmd_xbar_demux_001_src5_data                                                                      : std_logic_vector(75 downto 0); -- cmd_xbar_demux_001:src5_data -> pio_LEDR_s1_translator_avalon_universal_slave_0_agent:cp_data
	signal cmd_xbar_demux_001_src5_channel                                                                   : std_logic_vector(13 downto 0); -- cmd_xbar_demux_001:src5_channel -> pio_LEDR_s1_translator_avalon_universal_slave_0_agent:cp_channel
	signal cmd_xbar_demux_001_src6_endofpacket                                                               : std_logic;                     -- cmd_xbar_demux_001:src6_endofpacket -> pio_SW_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	signal cmd_xbar_demux_001_src6_valid                                                                     : std_logic;                     -- cmd_xbar_demux_001:src6_valid -> pio_SW_s1_translator_avalon_universal_slave_0_agent:cp_valid
	signal cmd_xbar_demux_001_src6_startofpacket                                                             : std_logic;                     -- cmd_xbar_demux_001:src6_startofpacket -> pio_SW_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	signal cmd_xbar_demux_001_src6_data                                                                      : std_logic_vector(75 downto 0); -- cmd_xbar_demux_001:src6_data -> pio_SW_s1_translator_avalon_universal_slave_0_agent:cp_data
	signal cmd_xbar_demux_001_src6_channel                                                                   : std_logic_vector(13 downto 0); -- cmd_xbar_demux_001:src6_channel -> pio_SW_s1_translator_avalon_universal_slave_0_agent:cp_channel
	signal cmd_xbar_demux_001_src7_endofpacket                                                               : std_logic;                     -- cmd_xbar_demux_001:src7_endofpacket -> pio_Button_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	signal cmd_xbar_demux_001_src7_valid                                                                     : std_logic;                     -- cmd_xbar_demux_001:src7_valid -> pio_Button_s1_translator_avalon_universal_slave_0_agent:cp_valid
	signal cmd_xbar_demux_001_src7_startofpacket                                                             : std_logic;                     -- cmd_xbar_demux_001:src7_startofpacket -> pio_Button_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	signal cmd_xbar_demux_001_src7_data                                                                      : std_logic_vector(75 downto 0); -- cmd_xbar_demux_001:src7_data -> pio_Button_s1_translator_avalon_universal_slave_0_agent:cp_data
	signal cmd_xbar_demux_001_src7_channel                                                                   : std_logic_vector(13 downto 0); -- cmd_xbar_demux_001:src7_channel -> pio_Button_s1_translator_avalon_universal_slave_0_agent:cp_channel
	signal cmd_xbar_demux_001_src8_endofpacket                                                               : std_logic;                     -- cmd_xbar_demux_001:src8_endofpacket -> lcd_control_slave_translator_avalon_universal_slave_0_agent:cp_endofpacket
	signal cmd_xbar_demux_001_src8_valid                                                                     : std_logic;                     -- cmd_xbar_demux_001:src8_valid -> lcd_control_slave_translator_avalon_universal_slave_0_agent:cp_valid
	signal cmd_xbar_demux_001_src8_startofpacket                                                             : std_logic;                     -- cmd_xbar_demux_001:src8_startofpacket -> lcd_control_slave_translator_avalon_universal_slave_0_agent:cp_startofpacket
	signal cmd_xbar_demux_001_src8_data                                                                      : std_logic_vector(75 downto 0); -- cmd_xbar_demux_001:src8_data -> lcd_control_slave_translator_avalon_universal_slave_0_agent:cp_data
	signal cmd_xbar_demux_001_src8_channel                                                                   : std_logic_vector(13 downto 0); -- cmd_xbar_demux_001:src8_channel -> lcd_control_slave_translator_avalon_universal_slave_0_agent:cp_channel
	signal cmd_xbar_demux_001_src9_endofpacket                                                               : std_logic;                     -- cmd_xbar_demux_001:src9_endofpacket -> uart_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	signal cmd_xbar_demux_001_src9_valid                                                                     : std_logic;                     -- cmd_xbar_demux_001:src9_valid -> uart_s1_translator_avalon_universal_slave_0_agent:cp_valid
	signal cmd_xbar_demux_001_src9_startofpacket                                                             : std_logic;                     -- cmd_xbar_demux_001:src9_startofpacket -> uart_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	signal cmd_xbar_demux_001_src9_data                                                                      : std_logic_vector(75 downto 0); -- cmd_xbar_demux_001:src9_data -> uart_s1_translator_avalon_universal_slave_0_agent:cp_data
	signal cmd_xbar_demux_001_src9_channel                                                                   : std_logic_vector(13 downto 0); -- cmd_xbar_demux_001:src9_channel -> uart_s1_translator_avalon_universal_slave_0_agent:cp_channel
	signal cmd_xbar_demux_001_src10_endofpacket                                                              : std_logic;                     -- cmd_xbar_demux_001:src10_endofpacket -> timer_0_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	signal cmd_xbar_demux_001_src10_valid                                                                    : std_logic;                     -- cmd_xbar_demux_001:src10_valid -> timer_0_s1_translator_avalon_universal_slave_0_agent:cp_valid
	signal cmd_xbar_demux_001_src10_startofpacket                                                            : std_logic;                     -- cmd_xbar_demux_001:src10_startofpacket -> timer_0_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	signal cmd_xbar_demux_001_src10_data                                                                     : std_logic_vector(75 downto 0); -- cmd_xbar_demux_001:src10_data -> timer_0_s1_translator_avalon_universal_slave_0_agent:cp_data
	signal cmd_xbar_demux_001_src10_channel                                                                  : std_logic_vector(13 downto 0); -- cmd_xbar_demux_001:src10_channel -> timer_0_s1_translator_avalon_universal_slave_0_agent:cp_channel
	signal cmd_xbar_demux_001_src11_endofpacket                                                              : std_logic;                     -- cmd_xbar_demux_001:src11_endofpacket -> pio_Data_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	signal cmd_xbar_demux_001_src11_valid                                                                    : std_logic;                     -- cmd_xbar_demux_001:src11_valid -> pio_Data_s1_translator_avalon_universal_slave_0_agent:cp_valid
	signal cmd_xbar_demux_001_src11_startofpacket                                                            : std_logic;                     -- cmd_xbar_demux_001:src11_startofpacket -> pio_Data_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	signal cmd_xbar_demux_001_src11_data                                                                     : std_logic_vector(75 downto 0); -- cmd_xbar_demux_001:src11_data -> pio_Data_s1_translator_avalon_universal_slave_0_agent:cp_data
	signal cmd_xbar_demux_001_src11_channel                                                                  : std_logic_vector(13 downto 0); -- cmd_xbar_demux_001:src11_channel -> pio_Data_s1_translator_avalon_universal_slave_0_agent:cp_channel
	signal cmd_xbar_demux_001_src12_endofpacket                                                              : std_logic;                     -- cmd_xbar_demux_001:src12_endofpacket -> pio_RdyData_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	signal cmd_xbar_demux_001_src12_valid                                                                    : std_logic;                     -- cmd_xbar_demux_001:src12_valid -> pio_RdyData_s1_translator_avalon_universal_slave_0_agent:cp_valid
	signal cmd_xbar_demux_001_src12_startofpacket                                                            : std_logic;                     -- cmd_xbar_demux_001:src12_startofpacket -> pio_RdyData_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	signal cmd_xbar_demux_001_src12_data                                                                     : std_logic_vector(75 downto 0); -- cmd_xbar_demux_001:src12_data -> pio_RdyData_s1_translator_avalon_universal_slave_0_agent:cp_data
	signal cmd_xbar_demux_001_src12_channel                                                                  : std_logic_vector(13 downto 0); -- cmd_xbar_demux_001:src12_channel -> pio_RdyData_s1_translator_avalon_universal_slave_0_agent:cp_channel
	signal cmd_xbar_demux_001_src13_endofpacket                                                              : std_logic;                     -- cmd_xbar_demux_001:src13_endofpacket -> pio_DataRead_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	signal cmd_xbar_demux_001_src13_valid                                                                    : std_logic;                     -- cmd_xbar_demux_001:src13_valid -> pio_DataRead_s1_translator_avalon_universal_slave_0_agent:cp_valid
	signal cmd_xbar_demux_001_src13_startofpacket                                                            : std_logic;                     -- cmd_xbar_demux_001:src13_startofpacket -> pio_DataRead_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	signal cmd_xbar_demux_001_src13_data                                                                     : std_logic_vector(75 downto 0); -- cmd_xbar_demux_001:src13_data -> pio_DataRead_s1_translator_avalon_universal_slave_0_agent:cp_data
	signal cmd_xbar_demux_001_src13_channel                                                                  : std_logic_vector(13 downto 0); -- cmd_xbar_demux_001:src13_channel -> pio_DataRead_s1_translator_avalon_universal_slave_0_agent:cp_channel
	signal rsp_xbar_demux_src0_endofpacket                                                                   : std_logic;                     -- rsp_xbar_demux:src0_endofpacket -> rsp_xbar_mux:sink0_endofpacket
	signal rsp_xbar_demux_src0_valid                                                                         : std_logic;                     -- rsp_xbar_demux:src0_valid -> rsp_xbar_mux:sink0_valid
	signal rsp_xbar_demux_src0_startofpacket                                                                 : std_logic;                     -- rsp_xbar_demux:src0_startofpacket -> rsp_xbar_mux:sink0_startofpacket
	signal rsp_xbar_demux_src0_data                                                                          : std_logic_vector(75 downto 0); -- rsp_xbar_demux:src0_data -> rsp_xbar_mux:sink0_data
	signal rsp_xbar_demux_src0_channel                                                                       : std_logic_vector(13 downto 0); -- rsp_xbar_demux:src0_channel -> rsp_xbar_mux:sink0_channel
	signal rsp_xbar_demux_src0_ready                                                                         : std_logic;                     -- rsp_xbar_mux:sink0_ready -> rsp_xbar_demux:src0_ready
	signal rsp_xbar_demux_src1_endofpacket                                                                   : std_logic;                     -- rsp_xbar_demux:src1_endofpacket -> rsp_xbar_mux_001:sink0_endofpacket
	signal rsp_xbar_demux_src1_valid                                                                         : std_logic;                     -- rsp_xbar_demux:src1_valid -> rsp_xbar_mux_001:sink0_valid
	signal rsp_xbar_demux_src1_startofpacket                                                                 : std_logic;                     -- rsp_xbar_demux:src1_startofpacket -> rsp_xbar_mux_001:sink0_startofpacket
	signal rsp_xbar_demux_src1_data                                                                          : std_logic_vector(75 downto 0); -- rsp_xbar_demux:src1_data -> rsp_xbar_mux_001:sink0_data
	signal rsp_xbar_demux_src1_channel                                                                       : std_logic_vector(13 downto 0); -- rsp_xbar_demux:src1_channel -> rsp_xbar_mux_001:sink0_channel
	signal rsp_xbar_demux_src1_ready                                                                         : std_logic;                     -- rsp_xbar_mux_001:sink0_ready -> rsp_xbar_demux:src1_ready
	signal rsp_xbar_demux_001_src0_endofpacket                                                               : std_logic;                     -- rsp_xbar_demux_001:src0_endofpacket -> rsp_xbar_mux:sink1_endofpacket
	signal rsp_xbar_demux_001_src0_valid                                                                     : std_logic;                     -- rsp_xbar_demux_001:src0_valid -> rsp_xbar_mux:sink1_valid
	signal rsp_xbar_demux_001_src0_startofpacket                                                             : std_logic;                     -- rsp_xbar_demux_001:src0_startofpacket -> rsp_xbar_mux:sink1_startofpacket
	signal rsp_xbar_demux_001_src0_data                                                                      : std_logic_vector(75 downto 0); -- rsp_xbar_demux_001:src0_data -> rsp_xbar_mux:sink1_data
	signal rsp_xbar_demux_001_src0_channel                                                                   : std_logic_vector(13 downto 0); -- rsp_xbar_demux_001:src0_channel -> rsp_xbar_mux:sink1_channel
	signal rsp_xbar_demux_001_src0_ready                                                                     : std_logic;                     -- rsp_xbar_mux:sink1_ready -> rsp_xbar_demux_001:src0_ready
	signal rsp_xbar_demux_001_src1_endofpacket                                                               : std_logic;                     -- rsp_xbar_demux_001:src1_endofpacket -> rsp_xbar_mux_001:sink1_endofpacket
	signal rsp_xbar_demux_001_src1_valid                                                                     : std_logic;                     -- rsp_xbar_demux_001:src1_valid -> rsp_xbar_mux_001:sink1_valid
	signal rsp_xbar_demux_001_src1_startofpacket                                                             : std_logic;                     -- rsp_xbar_demux_001:src1_startofpacket -> rsp_xbar_mux_001:sink1_startofpacket
	signal rsp_xbar_demux_001_src1_data                                                                      : std_logic_vector(75 downto 0); -- rsp_xbar_demux_001:src1_data -> rsp_xbar_mux_001:sink1_data
	signal rsp_xbar_demux_001_src1_channel                                                                   : std_logic_vector(13 downto 0); -- rsp_xbar_demux_001:src1_channel -> rsp_xbar_mux_001:sink1_channel
	signal rsp_xbar_demux_001_src1_ready                                                                     : std_logic;                     -- rsp_xbar_mux_001:sink1_ready -> rsp_xbar_demux_001:src1_ready
	signal rsp_xbar_demux_002_src0_endofpacket                                                               : std_logic;                     -- rsp_xbar_demux_002:src0_endofpacket -> rsp_xbar_mux_001:sink2_endofpacket
	signal rsp_xbar_demux_002_src0_valid                                                                     : std_logic;                     -- rsp_xbar_demux_002:src0_valid -> rsp_xbar_mux_001:sink2_valid
	signal rsp_xbar_demux_002_src0_startofpacket                                                             : std_logic;                     -- rsp_xbar_demux_002:src0_startofpacket -> rsp_xbar_mux_001:sink2_startofpacket
	signal rsp_xbar_demux_002_src0_data                                                                      : std_logic_vector(75 downto 0); -- rsp_xbar_demux_002:src0_data -> rsp_xbar_mux_001:sink2_data
	signal rsp_xbar_demux_002_src0_channel                                                                   : std_logic_vector(13 downto 0); -- rsp_xbar_demux_002:src0_channel -> rsp_xbar_mux_001:sink2_channel
	signal rsp_xbar_demux_002_src0_ready                                                                     : std_logic;                     -- rsp_xbar_mux_001:sink2_ready -> rsp_xbar_demux_002:src0_ready
	signal rsp_xbar_demux_003_src0_endofpacket                                                               : std_logic;                     -- rsp_xbar_demux_003:src0_endofpacket -> rsp_xbar_mux_001:sink3_endofpacket
	signal rsp_xbar_demux_003_src0_valid                                                                     : std_logic;                     -- rsp_xbar_demux_003:src0_valid -> rsp_xbar_mux_001:sink3_valid
	signal rsp_xbar_demux_003_src0_startofpacket                                                             : std_logic;                     -- rsp_xbar_demux_003:src0_startofpacket -> rsp_xbar_mux_001:sink3_startofpacket
	signal rsp_xbar_demux_003_src0_data                                                                      : std_logic_vector(75 downto 0); -- rsp_xbar_demux_003:src0_data -> rsp_xbar_mux_001:sink3_data
	signal rsp_xbar_demux_003_src0_channel                                                                   : std_logic_vector(13 downto 0); -- rsp_xbar_demux_003:src0_channel -> rsp_xbar_mux_001:sink3_channel
	signal rsp_xbar_demux_003_src0_ready                                                                     : std_logic;                     -- rsp_xbar_mux_001:sink3_ready -> rsp_xbar_demux_003:src0_ready
	signal rsp_xbar_demux_004_src0_endofpacket                                                               : std_logic;                     -- rsp_xbar_demux_004:src0_endofpacket -> rsp_xbar_mux_001:sink4_endofpacket
	signal rsp_xbar_demux_004_src0_valid                                                                     : std_logic;                     -- rsp_xbar_demux_004:src0_valid -> rsp_xbar_mux_001:sink4_valid
	signal rsp_xbar_demux_004_src0_startofpacket                                                             : std_logic;                     -- rsp_xbar_demux_004:src0_startofpacket -> rsp_xbar_mux_001:sink4_startofpacket
	signal rsp_xbar_demux_004_src0_data                                                                      : std_logic_vector(75 downto 0); -- rsp_xbar_demux_004:src0_data -> rsp_xbar_mux_001:sink4_data
	signal rsp_xbar_demux_004_src0_channel                                                                   : std_logic_vector(13 downto 0); -- rsp_xbar_demux_004:src0_channel -> rsp_xbar_mux_001:sink4_channel
	signal rsp_xbar_demux_004_src0_ready                                                                     : std_logic;                     -- rsp_xbar_mux_001:sink4_ready -> rsp_xbar_demux_004:src0_ready
	signal rsp_xbar_demux_005_src0_endofpacket                                                               : std_logic;                     -- rsp_xbar_demux_005:src0_endofpacket -> rsp_xbar_mux_001:sink5_endofpacket
	signal rsp_xbar_demux_005_src0_valid                                                                     : std_logic;                     -- rsp_xbar_demux_005:src0_valid -> rsp_xbar_mux_001:sink5_valid
	signal rsp_xbar_demux_005_src0_startofpacket                                                             : std_logic;                     -- rsp_xbar_demux_005:src0_startofpacket -> rsp_xbar_mux_001:sink5_startofpacket
	signal rsp_xbar_demux_005_src0_data                                                                      : std_logic_vector(75 downto 0); -- rsp_xbar_demux_005:src0_data -> rsp_xbar_mux_001:sink5_data
	signal rsp_xbar_demux_005_src0_channel                                                                   : std_logic_vector(13 downto 0); -- rsp_xbar_demux_005:src0_channel -> rsp_xbar_mux_001:sink5_channel
	signal rsp_xbar_demux_005_src0_ready                                                                     : std_logic;                     -- rsp_xbar_mux_001:sink5_ready -> rsp_xbar_demux_005:src0_ready
	signal rsp_xbar_demux_006_src0_endofpacket                                                               : std_logic;                     -- rsp_xbar_demux_006:src0_endofpacket -> rsp_xbar_mux_001:sink6_endofpacket
	signal rsp_xbar_demux_006_src0_valid                                                                     : std_logic;                     -- rsp_xbar_demux_006:src0_valid -> rsp_xbar_mux_001:sink6_valid
	signal rsp_xbar_demux_006_src0_startofpacket                                                             : std_logic;                     -- rsp_xbar_demux_006:src0_startofpacket -> rsp_xbar_mux_001:sink6_startofpacket
	signal rsp_xbar_demux_006_src0_data                                                                      : std_logic_vector(75 downto 0); -- rsp_xbar_demux_006:src0_data -> rsp_xbar_mux_001:sink6_data
	signal rsp_xbar_demux_006_src0_channel                                                                   : std_logic_vector(13 downto 0); -- rsp_xbar_demux_006:src0_channel -> rsp_xbar_mux_001:sink6_channel
	signal rsp_xbar_demux_006_src0_ready                                                                     : std_logic;                     -- rsp_xbar_mux_001:sink6_ready -> rsp_xbar_demux_006:src0_ready
	signal rsp_xbar_demux_007_src0_endofpacket                                                               : std_logic;                     -- rsp_xbar_demux_007:src0_endofpacket -> rsp_xbar_mux_001:sink7_endofpacket
	signal rsp_xbar_demux_007_src0_valid                                                                     : std_logic;                     -- rsp_xbar_demux_007:src0_valid -> rsp_xbar_mux_001:sink7_valid
	signal rsp_xbar_demux_007_src0_startofpacket                                                             : std_logic;                     -- rsp_xbar_demux_007:src0_startofpacket -> rsp_xbar_mux_001:sink7_startofpacket
	signal rsp_xbar_demux_007_src0_data                                                                      : std_logic_vector(75 downto 0); -- rsp_xbar_demux_007:src0_data -> rsp_xbar_mux_001:sink7_data
	signal rsp_xbar_demux_007_src0_channel                                                                   : std_logic_vector(13 downto 0); -- rsp_xbar_demux_007:src0_channel -> rsp_xbar_mux_001:sink7_channel
	signal rsp_xbar_demux_007_src0_ready                                                                     : std_logic;                     -- rsp_xbar_mux_001:sink7_ready -> rsp_xbar_demux_007:src0_ready
	signal rsp_xbar_demux_008_src0_endofpacket                                                               : std_logic;                     -- rsp_xbar_demux_008:src0_endofpacket -> rsp_xbar_mux_001:sink8_endofpacket
	signal rsp_xbar_demux_008_src0_valid                                                                     : std_logic;                     -- rsp_xbar_demux_008:src0_valid -> rsp_xbar_mux_001:sink8_valid
	signal rsp_xbar_demux_008_src0_startofpacket                                                             : std_logic;                     -- rsp_xbar_demux_008:src0_startofpacket -> rsp_xbar_mux_001:sink8_startofpacket
	signal rsp_xbar_demux_008_src0_data                                                                      : std_logic_vector(75 downto 0); -- rsp_xbar_demux_008:src0_data -> rsp_xbar_mux_001:sink8_data
	signal rsp_xbar_demux_008_src0_channel                                                                   : std_logic_vector(13 downto 0); -- rsp_xbar_demux_008:src0_channel -> rsp_xbar_mux_001:sink8_channel
	signal rsp_xbar_demux_008_src0_ready                                                                     : std_logic;                     -- rsp_xbar_mux_001:sink8_ready -> rsp_xbar_demux_008:src0_ready
	signal rsp_xbar_demux_009_src0_endofpacket                                                               : std_logic;                     -- rsp_xbar_demux_009:src0_endofpacket -> rsp_xbar_mux_001:sink9_endofpacket
	signal rsp_xbar_demux_009_src0_valid                                                                     : std_logic;                     -- rsp_xbar_demux_009:src0_valid -> rsp_xbar_mux_001:sink9_valid
	signal rsp_xbar_demux_009_src0_startofpacket                                                             : std_logic;                     -- rsp_xbar_demux_009:src0_startofpacket -> rsp_xbar_mux_001:sink9_startofpacket
	signal rsp_xbar_demux_009_src0_data                                                                      : std_logic_vector(75 downto 0); -- rsp_xbar_demux_009:src0_data -> rsp_xbar_mux_001:sink9_data
	signal rsp_xbar_demux_009_src0_channel                                                                   : std_logic_vector(13 downto 0); -- rsp_xbar_demux_009:src0_channel -> rsp_xbar_mux_001:sink9_channel
	signal rsp_xbar_demux_009_src0_ready                                                                     : std_logic;                     -- rsp_xbar_mux_001:sink9_ready -> rsp_xbar_demux_009:src0_ready
	signal rsp_xbar_demux_010_src0_endofpacket                                                               : std_logic;                     -- rsp_xbar_demux_010:src0_endofpacket -> rsp_xbar_mux_001:sink10_endofpacket
	signal rsp_xbar_demux_010_src0_valid                                                                     : std_logic;                     -- rsp_xbar_demux_010:src0_valid -> rsp_xbar_mux_001:sink10_valid
	signal rsp_xbar_demux_010_src0_startofpacket                                                             : std_logic;                     -- rsp_xbar_demux_010:src0_startofpacket -> rsp_xbar_mux_001:sink10_startofpacket
	signal rsp_xbar_demux_010_src0_data                                                                      : std_logic_vector(75 downto 0); -- rsp_xbar_demux_010:src0_data -> rsp_xbar_mux_001:sink10_data
	signal rsp_xbar_demux_010_src0_channel                                                                   : std_logic_vector(13 downto 0); -- rsp_xbar_demux_010:src0_channel -> rsp_xbar_mux_001:sink10_channel
	signal rsp_xbar_demux_010_src0_ready                                                                     : std_logic;                     -- rsp_xbar_mux_001:sink10_ready -> rsp_xbar_demux_010:src0_ready
	signal rsp_xbar_demux_011_src0_endofpacket                                                               : std_logic;                     -- rsp_xbar_demux_011:src0_endofpacket -> rsp_xbar_mux_001:sink11_endofpacket
	signal rsp_xbar_demux_011_src0_valid                                                                     : std_logic;                     -- rsp_xbar_demux_011:src0_valid -> rsp_xbar_mux_001:sink11_valid
	signal rsp_xbar_demux_011_src0_startofpacket                                                             : std_logic;                     -- rsp_xbar_demux_011:src0_startofpacket -> rsp_xbar_mux_001:sink11_startofpacket
	signal rsp_xbar_demux_011_src0_data                                                                      : std_logic_vector(75 downto 0); -- rsp_xbar_demux_011:src0_data -> rsp_xbar_mux_001:sink11_data
	signal rsp_xbar_demux_011_src0_channel                                                                   : std_logic_vector(13 downto 0); -- rsp_xbar_demux_011:src0_channel -> rsp_xbar_mux_001:sink11_channel
	signal rsp_xbar_demux_011_src0_ready                                                                     : std_logic;                     -- rsp_xbar_mux_001:sink11_ready -> rsp_xbar_demux_011:src0_ready
	signal rsp_xbar_demux_012_src0_endofpacket                                                               : std_logic;                     -- rsp_xbar_demux_012:src0_endofpacket -> rsp_xbar_mux_001:sink12_endofpacket
	signal rsp_xbar_demux_012_src0_valid                                                                     : std_logic;                     -- rsp_xbar_demux_012:src0_valid -> rsp_xbar_mux_001:sink12_valid
	signal rsp_xbar_demux_012_src0_startofpacket                                                             : std_logic;                     -- rsp_xbar_demux_012:src0_startofpacket -> rsp_xbar_mux_001:sink12_startofpacket
	signal rsp_xbar_demux_012_src0_data                                                                      : std_logic_vector(75 downto 0); -- rsp_xbar_demux_012:src0_data -> rsp_xbar_mux_001:sink12_data
	signal rsp_xbar_demux_012_src0_channel                                                                   : std_logic_vector(13 downto 0); -- rsp_xbar_demux_012:src0_channel -> rsp_xbar_mux_001:sink12_channel
	signal rsp_xbar_demux_012_src0_ready                                                                     : std_logic;                     -- rsp_xbar_mux_001:sink12_ready -> rsp_xbar_demux_012:src0_ready
	signal rsp_xbar_demux_013_src0_endofpacket                                                               : std_logic;                     -- rsp_xbar_demux_013:src0_endofpacket -> rsp_xbar_mux_001:sink13_endofpacket
	signal rsp_xbar_demux_013_src0_valid                                                                     : std_logic;                     -- rsp_xbar_demux_013:src0_valid -> rsp_xbar_mux_001:sink13_valid
	signal rsp_xbar_demux_013_src0_startofpacket                                                             : std_logic;                     -- rsp_xbar_demux_013:src0_startofpacket -> rsp_xbar_mux_001:sink13_startofpacket
	signal rsp_xbar_demux_013_src0_data                                                                      : std_logic_vector(75 downto 0); -- rsp_xbar_demux_013:src0_data -> rsp_xbar_mux_001:sink13_data
	signal rsp_xbar_demux_013_src0_channel                                                                   : std_logic_vector(13 downto 0); -- rsp_xbar_demux_013:src0_channel -> rsp_xbar_mux_001:sink13_channel
	signal rsp_xbar_demux_013_src0_ready                                                                     : std_logic;                     -- rsp_xbar_mux_001:sink13_ready -> rsp_xbar_demux_013:src0_ready
	signal limiter_cmd_src_endofpacket                                                                       : std_logic;                     -- limiter:cmd_src_endofpacket -> cmd_xbar_demux:sink_endofpacket
	signal limiter_cmd_src_startofpacket                                                                     : std_logic;                     -- limiter:cmd_src_startofpacket -> cmd_xbar_demux:sink_startofpacket
	signal limiter_cmd_src_data                                                                              : std_logic_vector(75 downto 0); -- limiter:cmd_src_data -> cmd_xbar_demux:sink_data
	signal limiter_cmd_src_channel                                                                           : std_logic_vector(13 downto 0); -- limiter:cmd_src_channel -> cmd_xbar_demux:sink_channel
	signal limiter_cmd_src_ready                                                                             : std_logic;                     -- cmd_xbar_demux:sink_ready -> limiter:cmd_src_ready
	signal rsp_xbar_mux_src_endofpacket                                                                      : std_logic;                     -- rsp_xbar_mux:src_endofpacket -> limiter:rsp_sink_endofpacket
	signal rsp_xbar_mux_src_valid                                                                            : std_logic;                     -- rsp_xbar_mux:src_valid -> limiter:rsp_sink_valid
	signal rsp_xbar_mux_src_startofpacket                                                                    : std_logic;                     -- rsp_xbar_mux:src_startofpacket -> limiter:rsp_sink_startofpacket
	signal rsp_xbar_mux_src_data                                                                             : std_logic_vector(75 downto 0); -- rsp_xbar_mux:src_data -> limiter:rsp_sink_data
	signal rsp_xbar_mux_src_channel                                                                          : std_logic_vector(13 downto 0); -- rsp_xbar_mux:src_channel -> limiter:rsp_sink_channel
	signal rsp_xbar_mux_src_ready                                                                            : std_logic;                     -- limiter:rsp_sink_ready -> rsp_xbar_mux:src_ready
	signal limiter_001_cmd_src_endofpacket                                                                   : std_logic;                     -- limiter_001:cmd_src_endofpacket -> cmd_xbar_demux_001:sink_endofpacket
	signal limiter_001_cmd_src_startofpacket                                                                 : std_logic;                     -- limiter_001:cmd_src_startofpacket -> cmd_xbar_demux_001:sink_startofpacket
	signal limiter_001_cmd_src_data                                                                          : std_logic_vector(75 downto 0); -- limiter_001:cmd_src_data -> cmd_xbar_demux_001:sink_data
	signal limiter_001_cmd_src_channel                                                                       : std_logic_vector(13 downto 0); -- limiter_001:cmd_src_channel -> cmd_xbar_demux_001:sink_channel
	signal limiter_001_cmd_src_ready                                                                         : std_logic;                     -- cmd_xbar_demux_001:sink_ready -> limiter_001:cmd_src_ready
	signal rsp_xbar_mux_001_src_endofpacket                                                                  : std_logic;                     -- rsp_xbar_mux_001:src_endofpacket -> limiter_001:rsp_sink_endofpacket
	signal rsp_xbar_mux_001_src_valid                                                                        : std_logic;                     -- rsp_xbar_mux_001:src_valid -> limiter_001:rsp_sink_valid
	signal rsp_xbar_mux_001_src_startofpacket                                                                : std_logic;                     -- rsp_xbar_mux_001:src_startofpacket -> limiter_001:rsp_sink_startofpacket
	signal rsp_xbar_mux_001_src_data                                                                         : std_logic_vector(75 downto 0); -- rsp_xbar_mux_001:src_data -> limiter_001:rsp_sink_data
	signal rsp_xbar_mux_001_src_channel                                                                      : std_logic_vector(13 downto 0); -- rsp_xbar_mux_001:src_channel -> limiter_001:rsp_sink_channel
	signal rsp_xbar_mux_001_src_ready                                                                        : std_logic;                     -- limiter_001:rsp_sink_ready -> rsp_xbar_mux_001:src_ready
	signal cmd_xbar_mux_src_endofpacket                                                                      : std_logic;                     -- cmd_xbar_mux:src_endofpacket -> nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent:cp_endofpacket
	signal cmd_xbar_mux_src_valid                                                                            : std_logic;                     -- cmd_xbar_mux:src_valid -> nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent:cp_valid
	signal cmd_xbar_mux_src_startofpacket                                                                    : std_logic;                     -- cmd_xbar_mux:src_startofpacket -> nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent:cp_startofpacket
	signal cmd_xbar_mux_src_data                                                                             : std_logic_vector(75 downto 0); -- cmd_xbar_mux:src_data -> nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent:cp_data
	signal cmd_xbar_mux_src_channel                                                                          : std_logic_vector(13 downto 0); -- cmd_xbar_mux:src_channel -> nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent:cp_channel
	signal cmd_xbar_mux_src_ready                                                                            : std_logic;                     -- nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_mux:src_ready
	signal id_router_src_endofpacket                                                                         : std_logic;                     -- id_router:src_endofpacket -> rsp_xbar_demux:sink_endofpacket
	signal id_router_src_valid                                                                               : std_logic;                     -- id_router:src_valid -> rsp_xbar_demux:sink_valid
	signal id_router_src_startofpacket                                                                       : std_logic;                     -- id_router:src_startofpacket -> rsp_xbar_demux:sink_startofpacket
	signal id_router_src_data                                                                                : std_logic_vector(75 downto 0); -- id_router:src_data -> rsp_xbar_demux:sink_data
	signal id_router_src_channel                                                                             : std_logic_vector(13 downto 0); -- id_router:src_channel -> rsp_xbar_demux:sink_channel
	signal id_router_src_ready                                                                               : std_logic;                     -- rsp_xbar_demux:sink_ready -> id_router:src_ready
	signal cmd_xbar_mux_001_src_endofpacket                                                                  : std_logic;                     -- cmd_xbar_mux_001:src_endofpacket -> onchip_memory_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	signal cmd_xbar_mux_001_src_valid                                                                        : std_logic;                     -- cmd_xbar_mux_001:src_valid -> onchip_memory_s1_translator_avalon_universal_slave_0_agent:cp_valid
	signal cmd_xbar_mux_001_src_startofpacket                                                                : std_logic;                     -- cmd_xbar_mux_001:src_startofpacket -> onchip_memory_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	signal cmd_xbar_mux_001_src_data                                                                         : std_logic_vector(75 downto 0); -- cmd_xbar_mux_001:src_data -> onchip_memory_s1_translator_avalon_universal_slave_0_agent:cp_data
	signal cmd_xbar_mux_001_src_channel                                                                      : std_logic_vector(13 downto 0); -- cmd_xbar_mux_001:src_channel -> onchip_memory_s1_translator_avalon_universal_slave_0_agent:cp_channel
	signal cmd_xbar_mux_001_src_ready                                                                        : std_logic;                     -- onchip_memory_s1_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_mux_001:src_ready
	signal id_router_001_src_endofpacket                                                                     : std_logic;                     -- id_router_001:src_endofpacket -> rsp_xbar_demux_001:sink_endofpacket
	signal id_router_001_src_valid                                                                           : std_logic;                     -- id_router_001:src_valid -> rsp_xbar_demux_001:sink_valid
	signal id_router_001_src_startofpacket                                                                   : std_logic;                     -- id_router_001:src_startofpacket -> rsp_xbar_demux_001:sink_startofpacket
	signal id_router_001_src_data                                                                            : std_logic_vector(75 downto 0); -- id_router_001:src_data -> rsp_xbar_demux_001:sink_data
	signal id_router_001_src_channel                                                                         : std_logic_vector(13 downto 0); -- id_router_001:src_channel -> rsp_xbar_demux_001:sink_channel
	signal id_router_001_src_ready                                                                           : std_logic;                     -- rsp_xbar_demux_001:sink_ready -> id_router_001:src_ready
	signal cmd_xbar_demux_001_src2_ready                                                                     : std_logic;                     -- jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_001:src2_ready
	signal id_router_002_src_endofpacket                                                                     : std_logic;                     -- id_router_002:src_endofpacket -> rsp_xbar_demux_002:sink_endofpacket
	signal id_router_002_src_valid                                                                           : std_logic;                     -- id_router_002:src_valid -> rsp_xbar_demux_002:sink_valid
	signal id_router_002_src_startofpacket                                                                   : std_logic;                     -- id_router_002:src_startofpacket -> rsp_xbar_demux_002:sink_startofpacket
	signal id_router_002_src_data                                                                            : std_logic_vector(75 downto 0); -- id_router_002:src_data -> rsp_xbar_demux_002:sink_data
	signal id_router_002_src_channel                                                                         : std_logic_vector(13 downto 0); -- id_router_002:src_channel -> rsp_xbar_demux_002:sink_channel
	signal id_router_002_src_ready                                                                           : std_logic;                     -- rsp_xbar_demux_002:sink_ready -> id_router_002:src_ready
	signal cmd_xbar_demux_001_src3_ready                                                                     : std_logic;                     -- sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_001:src3_ready
	signal id_router_003_src_endofpacket                                                                     : std_logic;                     -- id_router_003:src_endofpacket -> rsp_xbar_demux_003:sink_endofpacket
	signal id_router_003_src_valid                                                                           : std_logic;                     -- id_router_003:src_valid -> rsp_xbar_demux_003:sink_valid
	signal id_router_003_src_startofpacket                                                                   : std_logic;                     -- id_router_003:src_startofpacket -> rsp_xbar_demux_003:sink_startofpacket
	signal id_router_003_src_data                                                                            : std_logic_vector(75 downto 0); -- id_router_003:src_data -> rsp_xbar_demux_003:sink_data
	signal id_router_003_src_channel                                                                         : std_logic_vector(13 downto 0); -- id_router_003:src_channel -> rsp_xbar_demux_003:sink_channel
	signal id_router_003_src_ready                                                                           : std_logic;                     -- rsp_xbar_demux_003:sink_ready -> id_router_003:src_ready
	signal cmd_xbar_demux_001_src4_ready                                                                     : std_logic;                     -- pio_LEDG_s1_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_001:src4_ready
	signal id_router_004_src_endofpacket                                                                     : std_logic;                     -- id_router_004:src_endofpacket -> rsp_xbar_demux_004:sink_endofpacket
	signal id_router_004_src_valid                                                                           : std_logic;                     -- id_router_004:src_valid -> rsp_xbar_demux_004:sink_valid
	signal id_router_004_src_startofpacket                                                                   : std_logic;                     -- id_router_004:src_startofpacket -> rsp_xbar_demux_004:sink_startofpacket
	signal id_router_004_src_data                                                                            : std_logic_vector(75 downto 0); -- id_router_004:src_data -> rsp_xbar_demux_004:sink_data
	signal id_router_004_src_channel                                                                         : std_logic_vector(13 downto 0); -- id_router_004:src_channel -> rsp_xbar_demux_004:sink_channel
	signal id_router_004_src_ready                                                                           : std_logic;                     -- rsp_xbar_demux_004:sink_ready -> id_router_004:src_ready
	signal cmd_xbar_demux_001_src5_ready                                                                     : std_logic;                     -- pio_LEDR_s1_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_001:src5_ready
	signal id_router_005_src_endofpacket                                                                     : std_logic;                     -- id_router_005:src_endofpacket -> rsp_xbar_demux_005:sink_endofpacket
	signal id_router_005_src_valid                                                                           : std_logic;                     -- id_router_005:src_valid -> rsp_xbar_demux_005:sink_valid
	signal id_router_005_src_startofpacket                                                                   : std_logic;                     -- id_router_005:src_startofpacket -> rsp_xbar_demux_005:sink_startofpacket
	signal id_router_005_src_data                                                                            : std_logic_vector(75 downto 0); -- id_router_005:src_data -> rsp_xbar_demux_005:sink_data
	signal id_router_005_src_channel                                                                         : std_logic_vector(13 downto 0); -- id_router_005:src_channel -> rsp_xbar_demux_005:sink_channel
	signal id_router_005_src_ready                                                                           : std_logic;                     -- rsp_xbar_demux_005:sink_ready -> id_router_005:src_ready
	signal cmd_xbar_demux_001_src6_ready                                                                     : std_logic;                     -- pio_SW_s1_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_001:src6_ready
	signal id_router_006_src_endofpacket                                                                     : std_logic;                     -- id_router_006:src_endofpacket -> rsp_xbar_demux_006:sink_endofpacket
	signal id_router_006_src_valid                                                                           : std_logic;                     -- id_router_006:src_valid -> rsp_xbar_demux_006:sink_valid
	signal id_router_006_src_startofpacket                                                                   : std_logic;                     -- id_router_006:src_startofpacket -> rsp_xbar_demux_006:sink_startofpacket
	signal id_router_006_src_data                                                                            : std_logic_vector(75 downto 0); -- id_router_006:src_data -> rsp_xbar_demux_006:sink_data
	signal id_router_006_src_channel                                                                         : std_logic_vector(13 downto 0); -- id_router_006:src_channel -> rsp_xbar_demux_006:sink_channel
	signal id_router_006_src_ready                                                                           : std_logic;                     -- rsp_xbar_demux_006:sink_ready -> id_router_006:src_ready
	signal cmd_xbar_demux_001_src7_ready                                                                     : std_logic;                     -- pio_Button_s1_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_001:src7_ready
	signal id_router_007_src_endofpacket                                                                     : std_logic;                     -- id_router_007:src_endofpacket -> rsp_xbar_demux_007:sink_endofpacket
	signal id_router_007_src_valid                                                                           : std_logic;                     -- id_router_007:src_valid -> rsp_xbar_demux_007:sink_valid
	signal id_router_007_src_startofpacket                                                                   : std_logic;                     -- id_router_007:src_startofpacket -> rsp_xbar_demux_007:sink_startofpacket
	signal id_router_007_src_data                                                                            : std_logic_vector(75 downto 0); -- id_router_007:src_data -> rsp_xbar_demux_007:sink_data
	signal id_router_007_src_channel                                                                         : std_logic_vector(13 downto 0); -- id_router_007:src_channel -> rsp_xbar_demux_007:sink_channel
	signal id_router_007_src_ready                                                                           : std_logic;                     -- rsp_xbar_demux_007:sink_ready -> id_router_007:src_ready
	signal cmd_xbar_demux_001_src8_ready                                                                     : std_logic;                     -- lcd_control_slave_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_001:src8_ready
	signal id_router_008_src_endofpacket                                                                     : std_logic;                     -- id_router_008:src_endofpacket -> rsp_xbar_demux_008:sink_endofpacket
	signal id_router_008_src_valid                                                                           : std_logic;                     -- id_router_008:src_valid -> rsp_xbar_demux_008:sink_valid
	signal id_router_008_src_startofpacket                                                                   : std_logic;                     -- id_router_008:src_startofpacket -> rsp_xbar_demux_008:sink_startofpacket
	signal id_router_008_src_data                                                                            : std_logic_vector(75 downto 0); -- id_router_008:src_data -> rsp_xbar_demux_008:sink_data
	signal id_router_008_src_channel                                                                         : std_logic_vector(13 downto 0); -- id_router_008:src_channel -> rsp_xbar_demux_008:sink_channel
	signal id_router_008_src_ready                                                                           : std_logic;                     -- rsp_xbar_demux_008:sink_ready -> id_router_008:src_ready
	signal cmd_xbar_demux_001_src9_ready                                                                     : std_logic;                     -- uart_s1_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_001:src9_ready
	signal id_router_009_src_endofpacket                                                                     : std_logic;                     -- id_router_009:src_endofpacket -> rsp_xbar_demux_009:sink_endofpacket
	signal id_router_009_src_valid                                                                           : std_logic;                     -- id_router_009:src_valid -> rsp_xbar_demux_009:sink_valid
	signal id_router_009_src_startofpacket                                                                   : std_logic;                     -- id_router_009:src_startofpacket -> rsp_xbar_demux_009:sink_startofpacket
	signal id_router_009_src_data                                                                            : std_logic_vector(75 downto 0); -- id_router_009:src_data -> rsp_xbar_demux_009:sink_data
	signal id_router_009_src_channel                                                                         : std_logic_vector(13 downto 0); -- id_router_009:src_channel -> rsp_xbar_demux_009:sink_channel
	signal id_router_009_src_ready                                                                           : std_logic;                     -- rsp_xbar_demux_009:sink_ready -> id_router_009:src_ready
	signal cmd_xbar_demux_001_src10_ready                                                                    : std_logic;                     -- timer_0_s1_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_001:src10_ready
	signal id_router_010_src_endofpacket                                                                     : std_logic;                     -- id_router_010:src_endofpacket -> rsp_xbar_demux_010:sink_endofpacket
	signal id_router_010_src_valid                                                                           : std_logic;                     -- id_router_010:src_valid -> rsp_xbar_demux_010:sink_valid
	signal id_router_010_src_startofpacket                                                                   : std_logic;                     -- id_router_010:src_startofpacket -> rsp_xbar_demux_010:sink_startofpacket
	signal id_router_010_src_data                                                                            : std_logic_vector(75 downto 0); -- id_router_010:src_data -> rsp_xbar_demux_010:sink_data
	signal id_router_010_src_channel                                                                         : std_logic_vector(13 downto 0); -- id_router_010:src_channel -> rsp_xbar_demux_010:sink_channel
	signal id_router_010_src_ready                                                                           : std_logic;                     -- rsp_xbar_demux_010:sink_ready -> id_router_010:src_ready
	signal cmd_xbar_demux_001_src11_ready                                                                    : std_logic;                     -- pio_Data_s1_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_001:src11_ready
	signal id_router_011_src_endofpacket                                                                     : std_logic;                     -- id_router_011:src_endofpacket -> rsp_xbar_demux_011:sink_endofpacket
	signal id_router_011_src_valid                                                                           : std_logic;                     -- id_router_011:src_valid -> rsp_xbar_demux_011:sink_valid
	signal id_router_011_src_startofpacket                                                                   : std_logic;                     -- id_router_011:src_startofpacket -> rsp_xbar_demux_011:sink_startofpacket
	signal id_router_011_src_data                                                                            : std_logic_vector(75 downto 0); -- id_router_011:src_data -> rsp_xbar_demux_011:sink_data
	signal id_router_011_src_channel                                                                         : std_logic_vector(13 downto 0); -- id_router_011:src_channel -> rsp_xbar_demux_011:sink_channel
	signal id_router_011_src_ready                                                                           : std_logic;                     -- rsp_xbar_demux_011:sink_ready -> id_router_011:src_ready
	signal cmd_xbar_demux_001_src12_ready                                                                    : std_logic;                     -- pio_RdyData_s1_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_001:src12_ready
	signal id_router_012_src_endofpacket                                                                     : std_logic;                     -- id_router_012:src_endofpacket -> rsp_xbar_demux_012:sink_endofpacket
	signal id_router_012_src_valid                                                                           : std_logic;                     -- id_router_012:src_valid -> rsp_xbar_demux_012:sink_valid
	signal id_router_012_src_startofpacket                                                                   : std_logic;                     -- id_router_012:src_startofpacket -> rsp_xbar_demux_012:sink_startofpacket
	signal id_router_012_src_data                                                                            : std_logic_vector(75 downto 0); -- id_router_012:src_data -> rsp_xbar_demux_012:sink_data
	signal id_router_012_src_channel                                                                         : std_logic_vector(13 downto 0); -- id_router_012:src_channel -> rsp_xbar_demux_012:sink_channel
	signal id_router_012_src_ready                                                                           : std_logic;                     -- rsp_xbar_demux_012:sink_ready -> id_router_012:src_ready
	signal cmd_xbar_demux_001_src13_ready                                                                    : std_logic;                     -- pio_DataRead_s1_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_001:src13_ready
	signal id_router_013_src_endofpacket                                                                     : std_logic;                     -- id_router_013:src_endofpacket -> rsp_xbar_demux_013:sink_endofpacket
	signal id_router_013_src_valid                                                                           : std_logic;                     -- id_router_013:src_valid -> rsp_xbar_demux_013:sink_valid
	signal id_router_013_src_startofpacket                                                                   : std_logic;                     -- id_router_013:src_startofpacket -> rsp_xbar_demux_013:sink_startofpacket
	signal id_router_013_src_data                                                                            : std_logic_vector(75 downto 0); -- id_router_013:src_data -> rsp_xbar_demux_013:sink_data
	signal id_router_013_src_channel                                                                         : std_logic_vector(13 downto 0); -- id_router_013:src_channel -> rsp_xbar_demux_013:sink_channel
	signal id_router_013_src_ready                                                                           : std_logic;                     -- rsp_xbar_demux_013:sink_ready -> id_router_013:src_ready
	signal limiter_cmd_valid_data                                                                            : std_logic_vector(13 downto 0); -- limiter:cmd_src_valid -> cmd_xbar_demux:sink_valid
	signal limiter_001_cmd_valid_data                                                                        : std_logic_vector(13 downto 0); -- limiter_001:cmd_src_valid -> cmd_xbar_demux_001:sink_valid
	signal irq_mapper_receiver0_irq                                                                          : std_logic;                     -- jtag_uart:av_irq -> irq_mapper:receiver0_irq
	signal irq_mapper_receiver1_irq                                                                          : std_logic;                     -- timer_0:irq -> irq_mapper:receiver1_irq
	signal irq_mapper_receiver2_irq                                                                          : std_logic;                     -- uart:irq -> irq_mapper:receiver2_irq
	signal irq_mapper_receiver3_irq                                                                          : std_logic;                     -- pio_Button:irq -> irq_mapper:receiver3_irq
	signal irq_mapper_receiver4_irq                                                                          : std_logic;                     -- pio_RdyData:irq -> irq_mapper:receiver4_irq
	signal nios2_qsys_d_irq_irq                                                                              : std_logic_vector(31 downto 0); -- irq_mapper:sender_irq -> nios2_qsys:d_irq
	signal reset_reset_n_ports_inv                                                                           : std_logic;                     -- reset_reset_n:inv -> rst_controller:reset_in0
	signal jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_write_ports_inv                        : std_logic;                     -- jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_write:inv -> jtag_uart:av_write_n
	signal jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_read_ports_inv                         : std_logic;                     -- jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_read:inv -> jtag_uart:av_read_n
	signal pio_ledg_s1_translator_avalon_anti_slave_0_write_ports_inv                                        : std_logic;                     -- pio_ledg_s1_translator_avalon_anti_slave_0_write:inv -> pio_LEDG:write_n
	signal pio_ledr_s1_translator_avalon_anti_slave_0_write_ports_inv                                        : std_logic;                     -- pio_ledr_s1_translator_avalon_anti_slave_0_write:inv -> pio_LEDR:write_n
	signal pio_button_s1_translator_avalon_anti_slave_0_write_ports_inv                                      : std_logic;                     -- pio_button_s1_translator_avalon_anti_slave_0_write:inv -> pio_Button:write_n
	signal uart_s1_translator_avalon_anti_slave_0_write_ports_inv                                            : std_logic;                     -- uart_s1_translator_avalon_anti_slave_0_write:inv -> uart:write_n
	signal uart_s1_translator_avalon_anti_slave_0_read_ports_inv                                             : std_logic;                     -- uart_s1_translator_avalon_anti_slave_0_read:inv -> uart:read_n
	signal timer_0_s1_translator_avalon_anti_slave_0_write_ports_inv                                         : std_logic;                     -- timer_0_s1_translator_avalon_anti_slave_0_write:inv -> timer_0:write_n
	signal pio_rdydata_s1_translator_avalon_anti_slave_0_write_ports_inv                                     : std_logic;                     -- pio_rdydata_s1_translator_avalon_anti_slave_0_write:inv -> pio_RdyData:write_n
	signal pio_dataread_s1_translator_avalon_anti_slave_0_write_ports_inv                                    : std_logic;                     -- pio_dataread_s1_translator_avalon_anti_slave_0_write:inv -> pio_DataRead:write_n
	signal rst_controller_reset_out_reset_ports_inv                                                          : std_logic;                     -- rst_controller_reset_out_reset:inv -> [jtag_uart:rst_n, lcd:reset_n, nios2_qsys:reset_n, pio_Button:reset_n, pio_Data:reset_n, pio_DataRead:reset_n, pio_LEDG:reset_n, pio_LEDR:reset_n, pio_RdyData:reset_n, pio_SW:reset_n, sysid_qsys:reset_n, timer_0:reset_n, uart:reset_n]

begin

	nios2_qsys : component Nios1_nios2_qsys
		port map (
			clk                                   => clk_clk,                                                                   --                       clk.clk
			reset_n                               => rst_controller_reset_out_reset_ports_inv,                                  --                   reset_n.reset_n
			d_address                             => nios2_qsys_data_master_address,                                            --               data_master.address
			d_byteenable                          => nios2_qsys_data_master_byteenable,                                         --                          .byteenable
			d_read                                => nios2_qsys_data_master_read,                                               --                          .read
			d_readdata                            => nios2_qsys_data_master_readdata,                                           --                          .readdata
			d_waitrequest                         => nios2_qsys_data_master_waitrequest,                                        --                          .waitrequest
			d_write                               => nios2_qsys_data_master_write,                                              --                          .write
			d_writedata                           => nios2_qsys_data_master_writedata,                                          --                          .writedata
			d_readdatavalid                       => nios2_qsys_data_master_readdatavalid,                                      --                          .readdatavalid
			jtag_debug_module_debugaccess_to_roms => nios2_qsys_data_master_debugaccess,                                        --                          .debugaccess
			i_address                             => nios2_qsys_instruction_master_address,                                     --        instruction_master.address
			i_read                                => nios2_qsys_instruction_master_read,                                        --                          .read
			i_readdata                            => nios2_qsys_instruction_master_readdata,                                    --                          .readdata
			i_waitrequest                         => nios2_qsys_instruction_master_waitrequest,                                 --                          .waitrequest
			i_readdatavalid                       => nios2_qsys_instruction_master_readdatavalid,                               --                          .readdatavalid
			d_irq                                 => nios2_qsys_d_irq_irq,                                                      --                     d_irq.irq
			jtag_debug_module_resetrequest        => open,                                                                      --   jtag_debug_module_reset.reset
			jtag_debug_module_address             => nios2_qsys_jtag_debug_module_translator_avalon_anti_slave_0_address,       --         jtag_debug_module.address
			jtag_debug_module_begintransfer       => nios2_qsys_jtag_debug_module_translator_avalon_anti_slave_0_begintransfer, --                          .begintransfer
			jtag_debug_module_byteenable          => nios2_qsys_jtag_debug_module_translator_avalon_anti_slave_0_byteenable,    --                          .byteenable
			jtag_debug_module_debugaccess         => nios2_qsys_jtag_debug_module_translator_avalon_anti_slave_0_debugaccess,   --                          .debugaccess
			jtag_debug_module_readdata            => nios2_qsys_jtag_debug_module_translator_avalon_anti_slave_0_readdata,      --                          .readdata
			jtag_debug_module_select              => nios2_qsys_jtag_debug_module_translator_avalon_anti_slave_0_chipselect,    --                          .chipselect
			jtag_debug_module_write               => nios2_qsys_jtag_debug_module_translator_avalon_anti_slave_0_write,         --                          .write
			jtag_debug_module_writedata           => nios2_qsys_jtag_debug_module_translator_avalon_anti_slave_0_writedata,     --                          .writedata
			no_ci_readra                          => open                                                                       -- custom_instruction_master.readra
		);

	onchip_memory : component Nios1_onchip_memory
		port map (
			clk        => clk_clk,                                                    --   clk1.clk
			address    => onchip_memory_s1_translator_avalon_anti_slave_0_address,    --     s1.address
			chipselect => onchip_memory_s1_translator_avalon_anti_slave_0_chipselect, --       .chipselect
			clken      => onchip_memory_s1_translator_avalon_anti_slave_0_clken,      --       .clken
			readdata   => onchip_memory_s1_translator_avalon_anti_slave_0_readdata,   --       .readdata
			write      => onchip_memory_s1_translator_avalon_anti_slave_0_write,      --       .write
			writedata  => onchip_memory_s1_translator_avalon_anti_slave_0_writedata,  --       .writedata
			byteenable => onchip_memory_s1_translator_avalon_anti_slave_0_byteenable, --       .byteenable
			reset      => rst_controller_reset_out_reset                              -- reset1.reset
		);

	jtag_uart : component Nios1_jtag_uart
		port map (
			clk            => clk_clk,                                                                    --               clk.clk
			rst_n          => rst_controller_reset_out_reset_ports_inv,                                   --             reset.reset_n
			av_chipselect  => jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_chipselect,      -- avalon_jtag_slave.chipselect
			av_address     => jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_address,         --                  .address
			av_read_n      => jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_read_ports_inv,  --                  .read_n
			av_readdata    => jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_readdata,        --                  .readdata
			av_write_n     => jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_write_ports_inv, --                  .write_n
			av_writedata   => jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_writedata,       --                  .writedata
			av_waitrequest => jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_waitrequest,     --                  .waitrequest
			dataavailable  => open,                                                                       --                  .dataavailable
			readyfordata   => open,                                                                       --                  .readyfordata
			av_irq         => irq_mapper_receiver0_irq                                                    --               irq.irq
		);

	sysid_qsys : component Nios1_sysid_qsys
		port map (
			clock    => clk_clk,                                                          --           clk.clk
			reset_n  => rst_controller_reset_out_reset_ports_inv,                         --         reset.reset_n
			readdata => sysid_qsys_control_slave_translator_avalon_anti_slave_0_readdata, -- control_slave.readdata
			address  => sysid_qsys_control_slave_translator_avalon_anti_slave_0_address   --              .address
		);

	pio_ledg : component Nios1_pio_LEDG
		port map (
			clk        => clk_clk,                                                    --                 clk.clk
			reset_n    => rst_controller_reset_out_reset_ports_inv,                   --               reset.reset_n
			address    => pio_ledg_s1_translator_avalon_anti_slave_0_address,         --                  s1.address
			write_n    => pio_ledg_s1_translator_avalon_anti_slave_0_write_ports_inv, --                    .write_n
			writedata  => pio_ledg_s1_translator_avalon_anti_slave_0_writedata,       --                    .writedata
			chipselect => pio_ledg_s1_translator_avalon_anti_slave_0_chipselect,      --                    .chipselect
			readdata   => pio_ledg_s1_translator_avalon_anti_slave_0_readdata,        --                    .readdata
			out_port   => pio_ledg_export                                             -- external_connection.export
		);

	pio_ledr : component Nios1_pio_LEDR
		port map (
			clk        => clk_clk,                                                    --                 clk.clk
			reset_n    => rst_controller_reset_out_reset_ports_inv,                   --               reset.reset_n
			address    => pio_ledr_s1_translator_avalon_anti_slave_0_address,         --                  s1.address
			write_n    => pio_ledr_s1_translator_avalon_anti_slave_0_write_ports_inv, --                    .write_n
			writedata  => pio_ledr_s1_translator_avalon_anti_slave_0_writedata,       --                    .writedata
			chipselect => pio_ledr_s1_translator_avalon_anti_slave_0_chipselect,      --                    .chipselect
			readdata   => pio_ledr_s1_translator_avalon_anti_slave_0_readdata,        --                    .readdata
			out_port   => pio_ledr_export                                             -- external_connection.export
		);

	pio_sw : component Nios1_pio_SW
		port map (
			clk      => clk_clk,                                           --                 clk.clk
			reset_n  => rst_controller_reset_out_reset_ports_inv,          --               reset.reset_n
			address  => pio_sw_s1_translator_avalon_anti_slave_0_address,  --                  s1.address
			readdata => pio_sw_s1_translator_avalon_anti_slave_0_readdata, --                    .readdata
			in_port  => pio_sw_export                                      -- external_connection.export
		);

	pio_button : component Nios1_pio_Button
		port map (
			clk        => clk_clk,                                                      --                 clk.clk
			reset_n    => rst_controller_reset_out_reset_ports_inv,                     --               reset.reset_n
			address    => pio_button_s1_translator_avalon_anti_slave_0_address,         --                  s1.address
			write_n    => pio_button_s1_translator_avalon_anti_slave_0_write_ports_inv, --                    .write_n
			writedata  => pio_button_s1_translator_avalon_anti_slave_0_writedata,       --                    .writedata
			chipselect => pio_button_s1_translator_avalon_anti_slave_0_chipselect,      --                    .chipselect
			readdata   => pio_button_s1_translator_avalon_anti_slave_0_readdata,        --                    .readdata
			in_port    => pio_button_export,                                            -- external_connection.export
			irq        => irq_mapper_receiver3_irq                                      --                 irq.irq
		);

	lcd : component Nios1_lcd
		port map (
			clk           => clk_clk,                                                        --           clk.clk
			reset_n       => rst_controller_reset_out_reset_ports_inv,                       --         reset.reset_n
			address       => lcd_control_slave_translator_avalon_anti_slave_0_address,       -- control_slave.address
			begintransfer => lcd_control_slave_translator_avalon_anti_slave_0_begintransfer, --              .begintransfer
			read          => lcd_control_slave_translator_avalon_anti_slave_0_read,          --              .read
			readdata      => lcd_control_slave_translator_avalon_anti_slave_0_readdata,      --              .readdata
			write         => lcd_control_slave_translator_avalon_anti_slave_0_write,         --              .write
			writedata     => lcd_control_slave_translator_avalon_anti_slave_0_writedata,     --              .writedata
			LCD_data      => lcd_external_data,                                              --      external.export
			LCD_E         => lcd_external_E,                                                 --              .export
			LCD_RS        => lcd_external_RS,                                                --              .export
			LCD_RW        => lcd_external_RW                                                 --              .export
		);

	uart : component Nios1_uart
		port map (
			clk           => clk_clk,                                                --                 clk.clk
			reset_n       => rst_controller_reset_out_reset_ports_inv,               --               reset.reset_n
			address       => uart_s1_translator_avalon_anti_slave_0_address,         --                  s1.address
			begintransfer => uart_s1_translator_avalon_anti_slave_0_begintransfer,   --                    .begintransfer
			chipselect    => uart_s1_translator_avalon_anti_slave_0_chipselect,      --                    .chipselect
			read_n        => uart_s1_translator_avalon_anti_slave_0_read_ports_inv,  --                    .read_n
			write_n       => uart_s1_translator_avalon_anti_slave_0_write_ports_inv, --                    .write_n
			writedata     => uart_s1_translator_avalon_anti_slave_0_writedata,       --                    .writedata
			readdata      => uart_s1_translator_avalon_anti_slave_0_readdata,        --                    .readdata
			dataavailable => open,                                                   --                    .dataavailable
			readyfordata  => open,                                                   --                    .readyfordata
			rxd           => uart_external_rxd,                                      -- external_connection.export
			txd           => uart_external_txd,                                      --                    .export
			irq           => irq_mapper_receiver2_irq                                --                 irq.irq
		);

	timer_0 : component Nios1_timer_0
		port map (
			clk        => clk_clk,                                                   --   clk.clk
			reset_n    => rst_controller_reset_out_reset_ports_inv,                  -- reset.reset_n
			address    => timer_0_s1_translator_avalon_anti_slave_0_address,         --    s1.address
			writedata  => timer_0_s1_translator_avalon_anti_slave_0_writedata,       --      .writedata
			readdata   => timer_0_s1_translator_avalon_anti_slave_0_readdata,        --      .readdata
			chipselect => timer_0_s1_translator_avalon_anti_slave_0_chipselect,      --      .chipselect
			write_n    => timer_0_s1_translator_avalon_anti_slave_0_write_ports_inv, --      .write_n
			irq        => irq_mapper_receiver1_irq                                   --   irq.irq
		);

	pio_data : component Nios1_pio_Data
		port map (
			clk      => clk_clk,                                             --                 clk.clk
			reset_n  => rst_controller_reset_out_reset_ports_inv,            --               reset.reset_n
			address  => pio_data_s1_translator_avalon_anti_slave_0_address,  --                  s1.address
			readdata => pio_data_s1_translator_avalon_anti_slave_0_readdata, --                    .readdata
			in_port  => pio_data_export                                      -- external_connection.export
		);

	pio_rdydata : component Nios1_pio_RdyData
		port map (
			clk        => clk_clk,                                                       --                 clk.clk
			reset_n    => rst_controller_reset_out_reset_ports_inv,                      --               reset.reset_n
			address    => pio_rdydata_s1_translator_avalon_anti_slave_0_address,         --                  s1.address
			write_n    => pio_rdydata_s1_translator_avalon_anti_slave_0_write_ports_inv, --                    .write_n
			writedata  => pio_rdydata_s1_translator_avalon_anti_slave_0_writedata,       --                    .writedata
			chipselect => pio_rdydata_s1_translator_avalon_anti_slave_0_chipselect,      --                    .chipselect
			readdata   => pio_rdydata_s1_translator_avalon_anti_slave_0_readdata,        --                    .readdata
			in_port    => pio_rdydata_export,                                            -- external_connection.export
			irq        => irq_mapper_receiver4_irq                                       --                 irq.irq
		);

	pio_dataread : component Nios1_pio_DataRead
		port map (
			clk        => clk_clk,                                                        --                 clk.clk
			reset_n    => rst_controller_reset_out_reset_ports_inv,                       --               reset.reset_n
			address    => pio_dataread_s1_translator_avalon_anti_slave_0_address,         --                  s1.address
			write_n    => pio_dataread_s1_translator_avalon_anti_slave_0_write_ports_inv, --                    .write_n
			writedata  => pio_dataread_s1_translator_avalon_anti_slave_0_writedata,       --                    .writedata
			chipselect => pio_dataread_s1_translator_avalon_anti_slave_0_chipselect,      --                    .chipselect
			readdata   => pio_dataread_s1_translator_avalon_anti_slave_0_readdata,        --                    .readdata
			out_port   => pio_dataread_export                                             -- external_connection.export
		);

	nios2_qsys_instruction_master_translator : component Nios1_nios2_qsys_instruction_master_translator
		port map (
			clk               => clk_clk,                                                                          --                       clk.clk
			reset             => rst_controller_reset_out_reset,                                                   --                     reset.reset
			uav_address       => nios2_qsys_instruction_master_translator_avalon_universal_master_0_address,       -- avalon_universal_master_0.address
			uav_burstcount    => nios2_qsys_instruction_master_translator_avalon_universal_master_0_burstcount,    --                          .burstcount
			uav_read          => nios2_qsys_instruction_master_translator_avalon_universal_master_0_read,          --                          .read
			uav_write         => nios2_qsys_instruction_master_translator_avalon_universal_master_0_write,         --                          .write
			uav_waitrequest   => nios2_qsys_instruction_master_translator_avalon_universal_master_0_waitrequest,   --                          .waitrequest
			uav_readdatavalid => nios2_qsys_instruction_master_translator_avalon_universal_master_0_readdatavalid, --                          .readdatavalid
			uav_byteenable    => nios2_qsys_instruction_master_translator_avalon_universal_master_0_byteenable,    --                          .byteenable
			uav_readdata      => nios2_qsys_instruction_master_translator_avalon_universal_master_0_readdata,      --                          .readdata
			uav_writedata     => nios2_qsys_instruction_master_translator_avalon_universal_master_0_writedata,     --                          .writedata
			uav_lock          => nios2_qsys_instruction_master_translator_avalon_universal_master_0_lock,          --                          .lock
			uav_debugaccess   => nios2_qsys_instruction_master_translator_avalon_universal_master_0_debugaccess,   --                          .debugaccess
			av_address        => nios2_qsys_instruction_master_address,                                            --      avalon_anti_master_0.address
			av_waitrequest    => nios2_qsys_instruction_master_waitrequest,                                        --                          .waitrequest
			av_read           => nios2_qsys_instruction_master_read,                                               --                          .read
			av_readdata       => nios2_qsys_instruction_master_readdata,                                           --                          .readdata
			av_readdatavalid  => nios2_qsys_instruction_master_readdatavalid                                       --                          .readdatavalid
		);

	nios2_qsys_data_master_translator : component Nios1_nios2_qsys_data_master_translator
		port map (
			clk               => clk_clk,                                                                   --                       clk.clk
			reset             => rst_controller_reset_out_reset,                                            --                     reset.reset
			uav_address       => nios2_qsys_data_master_translator_avalon_universal_master_0_address,       -- avalon_universal_master_0.address
			uav_burstcount    => nios2_qsys_data_master_translator_avalon_universal_master_0_burstcount,    --                          .burstcount
			uav_read          => nios2_qsys_data_master_translator_avalon_universal_master_0_read,          --                          .read
			uav_write         => nios2_qsys_data_master_translator_avalon_universal_master_0_write,         --                          .write
			uav_waitrequest   => nios2_qsys_data_master_translator_avalon_universal_master_0_waitrequest,   --                          .waitrequest
			uav_readdatavalid => nios2_qsys_data_master_translator_avalon_universal_master_0_readdatavalid, --                          .readdatavalid
			uav_byteenable    => nios2_qsys_data_master_translator_avalon_universal_master_0_byteenable,    --                          .byteenable
			uav_readdata      => nios2_qsys_data_master_translator_avalon_universal_master_0_readdata,      --                          .readdata
			uav_writedata     => nios2_qsys_data_master_translator_avalon_universal_master_0_writedata,     --                          .writedata
			uav_lock          => nios2_qsys_data_master_translator_avalon_universal_master_0_lock,          --                          .lock
			uav_debugaccess   => nios2_qsys_data_master_translator_avalon_universal_master_0_debugaccess,   --                          .debugaccess
			av_address        => nios2_qsys_data_master_address,                                            --      avalon_anti_master_0.address
			av_waitrequest    => nios2_qsys_data_master_waitrequest,                                        --                          .waitrequest
			av_byteenable     => nios2_qsys_data_master_byteenable,                                         --                          .byteenable
			av_read           => nios2_qsys_data_master_read,                                               --                          .read
			av_readdata       => nios2_qsys_data_master_readdata,                                           --                          .readdata
			av_readdatavalid  => nios2_qsys_data_master_readdatavalid,                                      --                          .readdatavalid
			av_write          => nios2_qsys_data_master_write,                                              --                          .write
			av_writedata      => nios2_qsys_data_master_writedata,                                          --                          .writedata
			av_debugaccess    => nios2_qsys_data_master_debugaccess                                         --                          .debugaccess
		);

	nios2_qsys_jtag_debug_module_translator : component Nios1_nios2_qsys_jtag_debug_module_translator
		port map (
			clk               => clk_clk,                                                                                 --                      clk.clk
			reset             => rst_controller_reset_out_reset,                                                          --                    reset.reset
			uav_address       => nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_address,       -- avalon_universal_slave_0.address
			uav_burstcount    => nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_burstcount,    --                         .burstcount
			uav_read          => nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_read,          --                         .read
			uav_write         => nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_write,         --                         .write
			uav_waitrequest   => nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_waitrequest,   --                         .waitrequest
			uav_readdatavalid => nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_readdatavalid, --                         .readdatavalid
			uav_byteenable    => nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_byteenable,    --                         .byteenable
			uav_readdata      => nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_readdata,      --                         .readdata
			uav_writedata     => nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_writedata,     --                         .writedata
			uav_lock          => nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_lock,          --                         .lock
			uav_debugaccess   => nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_debugaccess,   --                         .debugaccess
			av_address        => nios2_qsys_jtag_debug_module_translator_avalon_anti_slave_0_address,                     --      avalon_anti_slave_0.address
			av_write          => nios2_qsys_jtag_debug_module_translator_avalon_anti_slave_0_write,                       --                         .write
			av_readdata       => nios2_qsys_jtag_debug_module_translator_avalon_anti_slave_0_readdata,                    --                         .readdata
			av_writedata      => nios2_qsys_jtag_debug_module_translator_avalon_anti_slave_0_writedata,                   --                         .writedata
			av_begintransfer  => nios2_qsys_jtag_debug_module_translator_avalon_anti_slave_0_begintransfer,               --                         .begintransfer
			av_byteenable     => nios2_qsys_jtag_debug_module_translator_avalon_anti_slave_0_byteenable,                  --                         .byteenable
			av_chipselect     => nios2_qsys_jtag_debug_module_translator_avalon_anti_slave_0_chipselect,                  --                         .chipselect
			av_debugaccess    => nios2_qsys_jtag_debug_module_translator_avalon_anti_slave_0_debugaccess                  --                         .debugaccess
		);

	onchip_memory_s1_translator : component Nios1_onchip_memory_s1_translator
		port map (
			clk               => clk_clk,                                                                     --                      clk.clk
			reset             => rst_controller_reset_out_reset,                                              --                    reset.reset
			uav_address       => onchip_memory_s1_translator_avalon_universal_slave_0_agent_m0_address,       -- avalon_universal_slave_0.address
			uav_burstcount    => onchip_memory_s1_translator_avalon_universal_slave_0_agent_m0_burstcount,    --                         .burstcount
			uav_read          => onchip_memory_s1_translator_avalon_universal_slave_0_agent_m0_read,          --                         .read
			uav_write         => onchip_memory_s1_translator_avalon_universal_slave_0_agent_m0_write,         --                         .write
			uav_waitrequest   => onchip_memory_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest,   --                         .waitrequest
			uav_readdatavalid => onchip_memory_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid, --                         .readdatavalid
			uav_byteenable    => onchip_memory_s1_translator_avalon_universal_slave_0_agent_m0_byteenable,    --                         .byteenable
			uav_readdata      => onchip_memory_s1_translator_avalon_universal_slave_0_agent_m0_readdata,      --                         .readdata
			uav_writedata     => onchip_memory_s1_translator_avalon_universal_slave_0_agent_m0_writedata,     --                         .writedata
			uav_lock          => onchip_memory_s1_translator_avalon_universal_slave_0_agent_m0_lock,          --                         .lock
			uav_debugaccess   => onchip_memory_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess,   --                         .debugaccess
			av_address        => onchip_memory_s1_translator_avalon_anti_slave_0_address,                     --      avalon_anti_slave_0.address
			av_write          => onchip_memory_s1_translator_avalon_anti_slave_0_write,                       --                         .write
			av_readdata       => onchip_memory_s1_translator_avalon_anti_slave_0_readdata,                    --                         .readdata
			av_writedata      => onchip_memory_s1_translator_avalon_anti_slave_0_writedata,                   --                         .writedata
			av_byteenable     => onchip_memory_s1_translator_avalon_anti_slave_0_byteenable,                  --                         .byteenable
			av_chipselect     => onchip_memory_s1_translator_avalon_anti_slave_0_chipselect,                  --                         .chipselect
			av_clken          => onchip_memory_s1_translator_avalon_anti_slave_0_clken                        --                         .clken
		);

	jtag_uart_avalon_jtag_slave_translator : component Nios1_jtag_uart_avalon_jtag_slave_translator
		port map (
			clk               => clk_clk,                                                                                --                      clk.clk
			reset             => rst_controller_reset_out_reset,                                                         --                    reset.reset
			uav_address       => jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_address,       -- avalon_universal_slave_0.address
			uav_burstcount    => jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_burstcount,    --                         .burstcount
			uav_read          => jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_read,          --                         .read
			uav_write         => jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_write,         --                         .write
			uav_waitrequest   => jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest,   --                         .waitrequest
			uav_readdatavalid => jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid, --                         .readdatavalid
			uav_byteenable    => jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_byteenable,    --                         .byteenable
			uav_readdata      => jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_readdata,      --                         .readdata
			uav_writedata     => jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_writedata,     --                         .writedata
			uav_lock          => jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_lock,          --                         .lock
			uav_debugaccess   => jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess,   --                         .debugaccess
			av_address        => jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_address,                     --      avalon_anti_slave_0.address
			av_write          => jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_write,                       --                         .write
			av_read           => jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_read,                        --                         .read
			av_readdata       => jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_readdata,                    --                         .readdata
			av_writedata      => jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_writedata,                   --                         .writedata
			av_waitrequest    => jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_waitrequest,                 --                         .waitrequest
			av_chipselect     => jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_chipselect                   --                         .chipselect
		);

	sysid_qsys_control_slave_translator : component Nios1_sysid_qsys_control_slave_translator
		port map (
			clk               => clk_clk,                                                                             --                      clk.clk
			reset             => rst_controller_reset_out_reset,                                                      --                    reset.reset
			uav_address       => sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent_m0_address,       -- avalon_universal_slave_0.address
			uav_burstcount    => sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent_m0_burstcount,    --                         .burstcount
			uav_read          => sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent_m0_read,          --                         .read
			uav_write         => sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent_m0_write,         --                         .write
			uav_waitrequest   => sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest,   --                         .waitrequest
			uav_readdatavalid => sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid, --                         .readdatavalid
			uav_byteenable    => sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent_m0_byteenable,    --                         .byteenable
			uav_readdata      => sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent_m0_readdata,      --                         .readdata
			uav_writedata     => sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent_m0_writedata,     --                         .writedata
			uav_lock          => sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent_m0_lock,          --                         .lock
			uav_debugaccess   => sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess,   --                         .debugaccess
			av_address        => sysid_qsys_control_slave_translator_avalon_anti_slave_0_address,                     --      avalon_anti_slave_0.address
			av_readdata       => sysid_qsys_control_slave_translator_avalon_anti_slave_0_readdata                     --                         .readdata
		);

	pio_ledg_s1_translator : component Nios1_pio_LEDG_s1_translator
		port map (
			clk               => clk_clk,                                                                --                      clk.clk
			reset             => rst_controller_reset_out_reset,                                         --                    reset.reset
			uav_address       => pio_ledg_s1_translator_avalon_universal_slave_0_agent_m0_address,       -- avalon_universal_slave_0.address
			uav_burstcount    => pio_ledg_s1_translator_avalon_universal_slave_0_agent_m0_burstcount,    --                         .burstcount
			uav_read          => pio_ledg_s1_translator_avalon_universal_slave_0_agent_m0_read,          --                         .read
			uav_write         => pio_ledg_s1_translator_avalon_universal_slave_0_agent_m0_write,         --                         .write
			uav_waitrequest   => pio_ledg_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest,   --                         .waitrequest
			uav_readdatavalid => pio_ledg_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid, --                         .readdatavalid
			uav_byteenable    => pio_ledg_s1_translator_avalon_universal_slave_0_agent_m0_byteenable,    --                         .byteenable
			uav_readdata      => pio_ledg_s1_translator_avalon_universal_slave_0_agent_m0_readdata,      --                         .readdata
			uav_writedata     => pio_ledg_s1_translator_avalon_universal_slave_0_agent_m0_writedata,     --                         .writedata
			uav_lock          => pio_ledg_s1_translator_avalon_universal_slave_0_agent_m0_lock,          --                         .lock
			uav_debugaccess   => pio_ledg_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess,   --                         .debugaccess
			av_address        => pio_ledg_s1_translator_avalon_anti_slave_0_address,                     --      avalon_anti_slave_0.address
			av_write          => pio_ledg_s1_translator_avalon_anti_slave_0_write,                       --                         .write
			av_readdata       => pio_ledg_s1_translator_avalon_anti_slave_0_readdata,                    --                         .readdata
			av_writedata      => pio_ledg_s1_translator_avalon_anti_slave_0_writedata,                   --                         .writedata
			av_chipselect     => pio_ledg_s1_translator_avalon_anti_slave_0_chipselect                   --                         .chipselect
		);

	pio_ledr_s1_translator : component Nios1_pio_LEDG_s1_translator
		port map (
			clk               => clk_clk,                                                                --                      clk.clk
			reset             => rst_controller_reset_out_reset,                                         --                    reset.reset
			uav_address       => pio_ledr_s1_translator_avalon_universal_slave_0_agent_m0_address,       -- avalon_universal_slave_0.address
			uav_burstcount    => pio_ledr_s1_translator_avalon_universal_slave_0_agent_m0_burstcount,    --                         .burstcount
			uav_read          => pio_ledr_s1_translator_avalon_universal_slave_0_agent_m0_read,          --                         .read
			uav_write         => pio_ledr_s1_translator_avalon_universal_slave_0_agent_m0_write,         --                         .write
			uav_waitrequest   => pio_ledr_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest,   --                         .waitrequest
			uav_readdatavalid => pio_ledr_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid, --                         .readdatavalid
			uav_byteenable    => pio_ledr_s1_translator_avalon_universal_slave_0_agent_m0_byteenable,    --                         .byteenable
			uav_readdata      => pio_ledr_s1_translator_avalon_universal_slave_0_agent_m0_readdata,      --                         .readdata
			uav_writedata     => pio_ledr_s1_translator_avalon_universal_slave_0_agent_m0_writedata,     --                         .writedata
			uav_lock          => pio_ledr_s1_translator_avalon_universal_slave_0_agent_m0_lock,          --                         .lock
			uav_debugaccess   => pio_ledr_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess,   --                         .debugaccess
			av_address        => pio_ledr_s1_translator_avalon_anti_slave_0_address,                     --      avalon_anti_slave_0.address
			av_write          => pio_ledr_s1_translator_avalon_anti_slave_0_write,                       --                         .write
			av_readdata       => pio_ledr_s1_translator_avalon_anti_slave_0_readdata,                    --                         .readdata
			av_writedata      => pio_ledr_s1_translator_avalon_anti_slave_0_writedata,                   --                         .writedata
			av_chipselect     => pio_ledr_s1_translator_avalon_anti_slave_0_chipselect                   --                         .chipselect
		);

	pio_sw_s1_translator : component Nios1_pio_SW_s1_translator
		port map (
			clk               => clk_clk,                                                              --                      clk.clk
			reset             => rst_controller_reset_out_reset,                                       --                    reset.reset
			uav_address       => pio_sw_s1_translator_avalon_universal_slave_0_agent_m0_address,       -- avalon_universal_slave_0.address
			uav_burstcount    => pio_sw_s1_translator_avalon_universal_slave_0_agent_m0_burstcount,    --                         .burstcount
			uav_read          => pio_sw_s1_translator_avalon_universal_slave_0_agent_m0_read,          --                         .read
			uav_write         => pio_sw_s1_translator_avalon_universal_slave_0_agent_m0_write,         --                         .write
			uav_waitrequest   => pio_sw_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest,   --                         .waitrequest
			uav_readdatavalid => pio_sw_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid, --                         .readdatavalid
			uav_byteenable    => pio_sw_s1_translator_avalon_universal_slave_0_agent_m0_byteenable,    --                         .byteenable
			uav_readdata      => pio_sw_s1_translator_avalon_universal_slave_0_agent_m0_readdata,      --                         .readdata
			uav_writedata     => pio_sw_s1_translator_avalon_universal_slave_0_agent_m0_writedata,     --                         .writedata
			uav_lock          => pio_sw_s1_translator_avalon_universal_slave_0_agent_m0_lock,          --                         .lock
			uav_debugaccess   => pio_sw_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess,   --                         .debugaccess
			av_address        => pio_sw_s1_translator_avalon_anti_slave_0_address,                     --      avalon_anti_slave_0.address
			av_readdata       => pio_sw_s1_translator_avalon_anti_slave_0_readdata                     --                         .readdata
		);

	pio_button_s1_translator : component Nios1_pio_Button_s1_translator
		port map (
			clk               => clk_clk,                                                                  --                      clk.clk
			reset             => rst_controller_reset_out_reset,                                           --                    reset.reset
			uav_address       => pio_button_s1_translator_avalon_universal_slave_0_agent_m0_address,       -- avalon_universal_slave_0.address
			uav_burstcount    => pio_button_s1_translator_avalon_universal_slave_0_agent_m0_burstcount,    --                         .burstcount
			uav_read          => pio_button_s1_translator_avalon_universal_slave_0_agent_m0_read,          --                         .read
			uav_write         => pio_button_s1_translator_avalon_universal_slave_0_agent_m0_write,         --                         .write
			uav_waitrequest   => pio_button_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest,   --                         .waitrequest
			uav_readdatavalid => pio_button_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid, --                         .readdatavalid
			uav_byteenable    => pio_button_s1_translator_avalon_universal_slave_0_agent_m0_byteenable,    --                         .byteenable
			uav_readdata      => pio_button_s1_translator_avalon_universal_slave_0_agent_m0_readdata,      --                         .readdata
			uav_writedata     => pio_button_s1_translator_avalon_universal_slave_0_agent_m0_writedata,     --                         .writedata
			uav_lock          => pio_button_s1_translator_avalon_universal_slave_0_agent_m0_lock,          --                         .lock
			uav_debugaccess   => pio_button_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess,   --                         .debugaccess
			av_address        => pio_button_s1_translator_avalon_anti_slave_0_address,                     --      avalon_anti_slave_0.address
			av_write          => pio_button_s1_translator_avalon_anti_slave_0_write,                       --                         .write
			av_readdata       => pio_button_s1_translator_avalon_anti_slave_0_readdata,                    --                         .readdata
			av_writedata      => pio_button_s1_translator_avalon_anti_slave_0_writedata,                   --                         .writedata
			av_chipselect     => pio_button_s1_translator_avalon_anti_slave_0_chipselect                   --                         .chipselect
		);

	lcd_control_slave_translator : component Nios1_lcd_control_slave_translator
		port map (
			clk               => clk_clk,                                                                      --                      clk.clk
			reset             => rst_controller_reset_out_reset,                                               --                    reset.reset
			uav_address       => lcd_control_slave_translator_avalon_universal_slave_0_agent_m0_address,       -- avalon_universal_slave_0.address
			uav_burstcount    => lcd_control_slave_translator_avalon_universal_slave_0_agent_m0_burstcount,    --                         .burstcount
			uav_read          => lcd_control_slave_translator_avalon_universal_slave_0_agent_m0_read,          --                         .read
			uav_write         => lcd_control_slave_translator_avalon_universal_slave_0_agent_m0_write,         --                         .write
			uav_waitrequest   => lcd_control_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest,   --                         .waitrequest
			uav_readdatavalid => lcd_control_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid, --                         .readdatavalid
			uav_byteenable    => lcd_control_slave_translator_avalon_universal_slave_0_agent_m0_byteenable,    --                         .byteenable
			uav_readdata      => lcd_control_slave_translator_avalon_universal_slave_0_agent_m0_readdata,      --                         .readdata
			uav_writedata     => lcd_control_slave_translator_avalon_universal_slave_0_agent_m0_writedata,     --                         .writedata
			uav_lock          => lcd_control_slave_translator_avalon_universal_slave_0_agent_m0_lock,          --                         .lock
			uav_debugaccess   => lcd_control_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess,   --                         .debugaccess
			av_address        => lcd_control_slave_translator_avalon_anti_slave_0_address,                     --      avalon_anti_slave_0.address
			av_write          => lcd_control_slave_translator_avalon_anti_slave_0_write,                       --                         .write
			av_read           => lcd_control_slave_translator_avalon_anti_slave_0_read,                        --                         .read
			av_readdata       => lcd_control_slave_translator_avalon_anti_slave_0_readdata,                    --                         .readdata
			av_writedata      => lcd_control_slave_translator_avalon_anti_slave_0_writedata,                   --                         .writedata
			av_begintransfer  => lcd_control_slave_translator_avalon_anti_slave_0_begintransfer                --                         .begintransfer
		);

	uart_s1_translator : component Nios1_uart_s1_translator
		port map (
			clk               => clk_clk,                                                            --                      clk.clk
			reset             => rst_controller_reset_out_reset,                                     --                    reset.reset
			uav_address       => uart_s1_translator_avalon_universal_slave_0_agent_m0_address,       -- avalon_universal_slave_0.address
			uav_burstcount    => uart_s1_translator_avalon_universal_slave_0_agent_m0_burstcount,    --                         .burstcount
			uav_read          => uart_s1_translator_avalon_universal_slave_0_agent_m0_read,          --                         .read
			uav_write         => uart_s1_translator_avalon_universal_slave_0_agent_m0_write,         --                         .write
			uav_waitrequest   => uart_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest,   --                         .waitrequest
			uav_readdatavalid => uart_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid, --                         .readdatavalid
			uav_byteenable    => uart_s1_translator_avalon_universal_slave_0_agent_m0_byteenable,    --                         .byteenable
			uav_readdata      => uart_s1_translator_avalon_universal_slave_0_agent_m0_readdata,      --                         .readdata
			uav_writedata     => uart_s1_translator_avalon_universal_slave_0_agent_m0_writedata,     --                         .writedata
			uav_lock          => uart_s1_translator_avalon_universal_slave_0_agent_m0_lock,          --                         .lock
			uav_debugaccess   => uart_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess,   --                         .debugaccess
			av_address        => uart_s1_translator_avalon_anti_slave_0_address,                     --      avalon_anti_slave_0.address
			av_write          => uart_s1_translator_avalon_anti_slave_0_write,                       --                         .write
			av_read           => uart_s1_translator_avalon_anti_slave_0_read,                        --                         .read
			av_readdata       => uart_s1_translator_avalon_anti_slave_0_readdata,                    --                         .readdata
			av_writedata      => uart_s1_translator_avalon_anti_slave_0_writedata,                   --                         .writedata
			av_begintransfer  => uart_s1_translator_avalon_anti_slave_0_begintransfer,               --                         .begintransfer
			av_chipselect     => uart_s1_translator_avalon_anti_slave_0_chipselect                   --                         .chipselect
		);

	timer_0_s1_translator : component Nios1_timer_0_s1_translator
		port map (
			clk               => clk_clk,                                                               --                      clk.clk
			reset             => rst_controller_reset_out_reset,                                        --                    reset.reset
			uav_address       => timer_0_s1_translator_avalon_universal_slave_0_agent_m0_address,       -- avalon_universal_slave_0.address
			uav_burstcount    => timer_0_s1_translator_avalon_universal_slave_0_agent_m0_burstcount,    --                         .burstcount
			uav_read          => timer_0_s1_translator_avalon_universal_slave_0_agent_m0_read,          --                         .read
			uav_write         => timer_0_s1_translator_avalon_universal_slave_0_agent_m0_write,         --                         .write
			uav_waitrequest   => timer_0_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest,   --                         .waitrequest
			uav_readdatavalid => timer_0_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid, --                         .readdatavalid
			uav_byteenable    => timer_0_s1_translator_avalon_universal_slave_0_agent_m0_byteenable,    --                         .byteenable
			uav_readdata      => timer_0_s1_translator_avalon_universal_slave_0_agent_m0_readdata,      --                         .readdata
			uav_writedata     => timer_0_s1_translator_avalon_universal_slave_0_agent_m0_writedata,     --                         .writedata
			uav_lock          => timer_0_s1_translator_avalon_universal_slave_0_agent_m0_lock,          --                         .lock
			uav_debugaccess   => timer_0_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess,   --                         .debugaccess
			av_address        => timer_0_s1_translator_avalon_anti_slave_0_address,                     --      avalon_anti_slave_0.address
			av_write          => timer_0_s1_translator_avalon_anti_slave_0_write,                       --                         .write
			av_readdata       => timer_0_s1_translator_avalon_anti_slave_0_readdata,                    --                         .readdata
			av_writedata      => timer_0_s1_translator_avalon_anti_slave_0_writedata,                   --                         .writedata
			av_chipselect     => timer_0_s1_translator_avalon_anti_slave_0_chipselect                   --                         .chipselect
		);

	pio_data_s1_translator : component Nios1_pio_SW_s1_translator
		port map (
			clk               => clk_clk,                                                                --                      clk.clk
			reset             => rst_controller_reset_out_reset,                                         --                    reset.reset
			uav_address       => pio_data_s1_translator_avalon_universal_slave_0_agent_m0_address,       -- avalon_universal_slave_0.address
			uav_burstcount    => pio_data_s1_translator_avalon_universal_slave_0_agent_m0_burstcount,    --                         .burstcount
			uav_read          => pio_data_s1_translator_avalon_universal_slave_0_agent_m0_read,          --                         .read
			uav_write         => pio_data_s1_translator_avalon_universal_slave_0_agent_m0_write,         --                         .write
			uav_waitrequest   => pio_data_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest,   --                         .waitrequest
			uav_readdatavalid => pio_data_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid, --                         .readdatavalid
			uav_byteenable    => pio_data_s1_translator_avalon_universal_slave_0_agent_m0_byteenable,    --                         .byteenable
			uav_readdata      => pio_data_s1_translator_avalon_universal_slave_0_agent_m0_readdata,      --                         .readdata
			uav_writedata     => pio_data_s1_translator_avalon_universal_slave_0_agent_m0_writedata,     --                         .writedata
			uav_lock          => pio_data_s1_translator_avalon_universal_slave_0_agent_m0_lock,          --                         .lock
			uav_debugaccess   => pio_data_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess,   --                         .debugaccess
			av_address        => pio_data_s1_translator_avalon_anti_slave_0_address,                     --      avalon_anti_slave_0.address
			av_readdata       => pio_data_s1_translator_avalon_anti_slave_0_readdata                     --                         .readdata
		);

	pio_rdydata_s1_translator : component Nios1_pio_Button_s1_translator
		port map (
			clk               => clk_clk,                                                                   --                      clk.clk
			reset             => rst_controller_reset_out_reset,                                            --                    reset.reset
			uav_address       => pio_rdydata_s1_translator_avalon_universal_slave_0_agent_m0_address,       -- avalon_universal_slave_0.address
			uav_burstcount    => pio_rdydata_s1_translator_avalon_universal_slave_0_agent_m0_burstcount,    --                         .burstcount
			uav_read          => pio_rdydata_s1_translator_avalon_universal_slave_0_agent_m0_read,          --                         .read
			uav_write         => pio_rdydata_s1_translator_avalon_universal_slave_0_agent_m0_write,         --                         .write
			uav_waitrequest   => pio_rdydata_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest,   --                         .waitrequest
			uav_readdatavalid => pio_rdydata_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid, --                         .readdatavalid
			uav_byteenable    => pio_rdydata_s1_translator_avalon_universal_slave_0_agent_m0_byteenable,    --                         .byteenable
			uav_readdata      => pio_rdydata_s1_translator_avalon_universal_slave_0_agent_m0_readdata,      --                         .readdata
			uav_writedata     => pio_rdydata_s1_translator_avalon_universal_slave_0_agent_m0_writedata,     --                         .writedata
			uav_lock          => pio_rdydata_s1_translator_avalon_universal_slave_0_agent_m0_lock,          --                         .lock
			uav_debugaccess   => pio_rdydata_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess,   --                         .debugaccess
			av_address        => pio_rdydata_s1_translator_avalon_anti_slave_0_address,                     --      avalon_anti_slave_0.address
			av_write          => pio_rdydata_s1_translator_avalon_anti_slave_0_write,                       --                         .write
			av_readdata       => pio_rdydata_s1_translator_avalon_anti_slave_0_readdata,                    --                         .readdata
			av_writedata      => pio_rdydata_s1_translator_avalon_anti_slave_0_writedata,                   --                         .writedata
			av_chipselect     => pio_rdydata_s1_translator_avalon_anti_slave_0_chipselect                   --                         .chipselect
		);

	pio_dataread_s1_translator : component Nios1_pio_LEDG_s1_translator
		port map (
			clk               => clk_clk,                                                                    --                      clk.clk
			reset             => rst_controller_reset_out_reset,                                             --                    reset.reset
			uav_address       => pio_dataread_s1_translator_avalon_universal_slave_0_agent_m0_address,       -- avalon_universal_slave_0.address
			uav_burstcount    => pio_dataread_s1_translator_avalon_universal_slave_0_agent_m0_burstcount,    --                         .burstcount
			uav_read          => pio_dataread_s1_translator_avalon_universal_slave_0_agent_m0_read,          --                         .read
			uav_write         => pio_dataread_s1_translator_avalon_universal_slave_0_agent_m0_write,         --                         .write
			uav_waitrequest   => pio_dataread_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest,   --                         .waitrequest
			uav_readdatavalid => pio_dataread_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid, --                         .readdatavalid
			uav_byteenable    => pio_dataread_s1_translator_avalon_universal_slave_0_agent_m0_byteenable,    --                         .byteenable
			uav_readdata      => pio_dataread_s1_translator_avalon_universal_slave_0_agent_m0_readdata,      --                         .readdata
			uav_writedata     => pio_dataread_s1_translator_avalon_universal_slave_0_agent_m0_writedata,     --                         .writedata
			uav_lock          => pio_dataread_s1_translator_avalon_universal_slave_0_agent_m0_lock,          --                         .lock
			uav_debugaccess   => pio_dataread_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess,   --                         .debugaccess
			av_address        => pio_dataread_s1_translator_avalon_anti_slave_0_address,                     --      avalon_anti_slave_0.address
			av_write          => pio_dataread_s1_translator_avalon_anti_slave_0_write,                       --                         .write
			av_readdata       => pio_dataread_s1_translator_avalon_anti_slave_0_readdata,                    --                         .readdata
			av_writedata      => pio_dataread_s1_translator_avalon_anti_slave_0_writedata,                   --                         .writedata
			av_chipselect     => pio_dataread_s1_translator_avalon_anti_slave_0_chipselect                   --                         .chipselect
		);

	pio_ledg_s1_translator_avalon_universal_slave_0_agent : component Nios1_pio_LEDG_s1_translator_avalon_universal_slave_0_agent
		port map (
			clk                     => clk_clk,                                                                          --             clk.clk
			reset                   => rst_controller_reset_out_reset,                                                   --       clk_reset.reset
			m0_address              => pio_ledg_s1_translator_avalon_universal_slave_0_agent_m0_address,                 --              m0.address
			m0_burstcount           => pio_ledg_s1_translator_avalon_universal_slave_0_agent_m0_burstcount,              --                .burstcount
			m0_byteenable           => pio_ledg_s1_translator_avalon_universal_slave_0_agent_m0_byteenable,              --                .byteenable
			m0_debugaccess          => pio_ledg_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess,             --                .debugaccess
			m0_lock                 => pio_ledg_s1_translator_avalon_universal_slave_0_agent_m0_lock,                    --                .lock
			m0_readdata             => pio_ledg_s1_translator_avalon_universal_slave_0_agent_m0_readdata,                --                .readdata
			m0_readdatavalid        => pio_ledg_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid,           --                .readdatavalid
			m0_read                 => pio_ledg_s1_translator_avalon_universal_slave_0_agent_m0_read,                    --                .read
			m0_waitrequest          => pio_ledg_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest,             --                .waitrequest
			m0_writedata            => pio_ledg_s1_translator_avalon_universal_slave_0_agent_m0_writedata,               --                .writedata
			m0_write                => pio_ledg_s1_translator_avalon_universal_slave_0_agent_m0_write,                   --                .write
			rp_endofpacket          => pio_ledg_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket,             --              rp.endofpacket
			rp_ready                => pio_ledg_s1_translator_avalon_universal_slave_0_agent_rp_ready,                   --                .ready
			rp_valid                => pio_ledg_s1_translator_avalon_universal_slave_0_agent_rp_valid,                   --                .valid
			rp_data                 => pio_ledg_s1_translator_avalon_universal_slave_0_agent_rp_data,                    --                .data
			rp_startofpacket        => pio_ledg_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket,           --                .startofpacket
			cp_ready                => cmd_xbar_demux_001_src4_ready,                                                    --              cp.ready
			cp_valid                => cmd_xbar_demux_001_src4_valid,                                                    --                .valid
			cp_data                 => cmd_xbar_demux_001_src4_data,                                                     --                .data
			cp_startofpacket        => cmd_xbar_demux_001_src4_startofpacket,                                            --                .startofpacket
			cp_endofpacket          => cmd_xbar_demux_001_src4_endofpacket,                                              --                .endofpacket
			cp_channel              => cmd_xbar_demux_001_src4_channel,                                                  --                .channel
			rf_sink_ready           => pio_ledg_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready,         --         rf_sink.ready
			rf_sink_valid           => pio_ledg_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid,         --                .valid
			rf_sink_startofpacket   => pio_ledg_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket, --                .startofpacket
			rf_sink_endofpacket     => pio_ledg_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket,   --                .endofpacket
			rf_sink_data            => pio_ledg_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data,          --                .data
			rf_source_ready         => pio_ledg_s1_translator_avalon_universal_slave_0_agent_rf_source_ready,            --       rf_source.ready
			rf_source_valid         => pio_ledg_s1_translator_avalon_universal_slave_0_agent_rf_source_valid,            --                .valid
			rf_source_startofpacket => pio_ledg_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket,    --                .startofpacket
			rf_source_endofpacket   => pio_ledg_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket,      --                .endofpacket
			rf_source_data          => pio_ledg_s1_translator_avalon_universal_slave_0_agent_rf_source_data,             --                .data
			rdata_fifo_sink_ready   => pio_ledg_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready,       -- rdata_fifo_sink.ready
			rdata_fifo_sink_valid   => pio_ledg_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid,       --                .valid
			rdata_fifo_sink_data    => pio_ledg_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data,        --                .data
			rdata_fifo_src_ready    => pio_ledg_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready,       --  rdata_fifo_src.ready
			rdata_fifo_src_valid    => pio_ledg_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid,       --                .valid
			rdata_fifo_src_data     => pio_ledg_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data         --                .data
		);

	pio_ledg_s1_translator_avalon_universal_slave_0_agent_rsp_fifo : component Nios1_pio_LEDG_s1_translator_avalon_universal_slave_0_agent_rsp_fifo
		port map (
			clk               => clk_clk,                                                                          --       clk.clk
			reset             => rst_controller_reset_out_reset,                                                   -- clk_reset.reset
			in_data           => pio_ledg_s1_translator_avalon_universal_slave_0_agent_rf_source_data,             --        in.data
			in_valid          => pio_ledg_s1_translator_avalon_universal_slave_0_agent_rf_source_valid,            --          .valid
			in_ready          => pio_ledg_s1_translator_avalon_universal_slave_0_agent_rf_source_ready,            --          .ready
			in_startofpacket  => pio_ledg_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket,    --          .startofpacket
			in_endofpacket    => pio_ledg_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket,      --          .endofpacket
			out_data          => pio_ledg_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data,          --       out.data
			out_valid         => pio_ledg_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid,         --          .valid
			out_ready         => pio_ledg_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready,         --          .ready
			out_startofpacket => pio_ledg_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket, --          .startofpacket
			out_endofpacket   => pio_ledg_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket    --          .endofpacket
		);

	pio_ledr_s1_translator_avalon_universal_slave_0_agent : component Nios1_pio_LEDR_s1_translator_avalon_universal_slave_0_agent
		port map (
			clk                     => clk_clk,                                                                          --             clk.clk
			reset                   => rst_controller_reset_out_reset,                                                   --       clk_reset.reset
			m0_address              => pio_ledr_s1_translator_avalon_universal_slave_0_agent_m0_address,                 --              m0.address
			m0_burstcount           => pio_ledr_s1_translator_avalon_universal_slave_0_agent_m0_burstcount,              --                .burstcount
			m0_byteenable           => pio_ledr_s1_translator_avalon_universal_slave_0_agent_m0_byteenable,              --                .byteenable
			m0_debugaccess          => pio_ledr_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess,             --                .debugaccess
			m0_lock                 => pio_ledr_s1_translator_avalon_universal_slave_0_agent_m0_lock,                    --                .lock
			m0_readdata             => pio_ledr_s1_translator_avalon_universal_slave_0_agent_m0_readdata,                --                .readdata
			m0_readdatavalid        => pio_ledr_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid,           --                .readdatavalid
			m0_read                 => pio_ledr_s1_translator_avalon_universal_slave_0_agent_m0_read,                    --                .read
			m0_waitrequest          => pio_ledr_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest,             --                .waitrequest
			m0_writedata            => pio_ledr_s1_translator_avalon_universal_slave_0_agent_m0_writedata,               --                .writedata
			m0_write                => pio_ledr_s1_translator_avalon_universal_slave_0_agent_m0_write,                   --                .write
			rp_endofpacket          => pio_ledr_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket,             --              rp.endofpacket
			rp_ready                => pio_ledr_s1_translator_avalon_universal_slave_0_agent_rp_ready,                   --                .ready
			rp_valid                => pio_ledr_s1_translator_avalon_universal_slave_0_agent_rp_valid,                   --                .valid
			rp_data                 => pio_ledr_s1_translator_avalon_universal_slave_0_agent_rp_data,                    --                .data
			rp_startofpacket        => pio_ledr_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket,           --                .startofpacket
			cp_ready                => cmd_xbar_demux_001_src5_ready,                                                    --              cp.ready
			cp_valid                => cmd_xbar_demux_001_src5_valid,                                                    --                .valid
			cp_data                 => cmd_xbar_demux_001_src5_data,                                                     --                .data
			cp_startofpacket        => cmd_xbar_demux_001_src5_startofpacket,                                            --                .startofpacket
			cp_endofpacket          => cmd_xbar_demux_001_src5_endofpacket,                                              --                .endofpacket
			cp_channel              => cmd_xbar_demux_001_src5_channel,                                                  --                .channel
			rf_sink_ready           => pio_ledr_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready,         --         rf_sink.ready
			rf_sink_valid           => pio_ledr_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid,         --                .valid
			rf_sink_startofpacket   => pio_ledr_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket, --                .startofpacket
			rf_sink_endofpacket     => pio_ledr_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket,   --                .endofpacket
			rf_sink_data            => pio_ledr_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data,          --                .data
			rf_source_ready         => pio_ledr_s1_translator_avalon_universal_slave_0_agent_rf_source_ready,            --       rf_source.ready
			rf_source_valid         => pio_ledr_s1_translator_avalon_universal_slave_0_agent_rf_source_valid,            --                .valid
			rf_source_startofpacket => pio_ledr_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket,    --                .startofpacket
			rf_source_endofpacket   => pio_ledr_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket,      --                .endofpacket
			rf_source_data          => pio_ledr_s1_translator_avalon_universal_slave_0_agent_rf_source_data,             --                .data
			rdata_fifo_sink_ready   => pio_ledr_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready,       -- rdata_fifo_sink.ready
			rdata_fifo_sink_valid   => pio_ledr_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid,       --                .valid
			rdata_fifo_sink_data    => pio_ledr_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data,        --                .data
			rdata_fifo_src_ready    => pio_ledr_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready,       --  rdata_fifo_src.ready
			rdata_fifo_src_valid    => pio_ledr_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid,       --                .valid
			rdata_fifo_src_data     => pio_ledr_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data         --                .data
		);

	pio_ledr_s1_translator_avalon_universal_slave_0_agent_rsp_fifo : component Nios1_pio_LEDG_s1_translator_avalon_universal_slave_0_agent_rsp_fifo
		port map (
			clk               => clk_clk,                                                                          --       clk.clk
			reset             => rst_controller_reset_out_reset,                                                   -- clk_reset.reset
			in_data           => pio_ledr_s1_translator_avalon_universal_slave_0_agent_rf_source_data,             --        in.data
			in_valid          => pio_ledr_s1_translator_avalon_universal_slave_0_agent_rf_source_valid,            --          .valid
			in_ready          => pio_ledr_s1_translator_avalon_universal_slave_0_agent_rf_source_ready,            --          .ready
			in_startofpacket  => pio_ledr_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket,    --          .startofpacket
			in_endofpacket    => pio_ledr_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket,      --          .endofpacket
			out_data          => pio_ledr_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data,          --       out.data
			out_valid         => pio_ledr_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid,         --          .valid
			out_ready         => pio_ledr_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready,         --          .ready
			out_startofpacket => pio_ledr_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket, --          .startofpacket
			out_endofpacket   => pio_ledr_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket    --          .endofpacket
		);

	sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent : component Nios1_sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent
		port map (
			clk                     => clk_clk,                                                                                       --             clk.clk
			reset                   => rst_controller_reset_out_reset,                                                                --       clk_reset.reset
			m0_address              => sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent_m0_address,                 --              m0.address
			m0_burstcount           => sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent_m0_burstcount,              --                .burstcount
			m0_byteenable           => sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent_m0_byteenable,              --                .byteenable
			m0_debugaccess          => sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess,             --                .debugaccess
			m0_lock                 => sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent_m0_lock,                    --                .lock
			m0_readdata             => sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent_m0_readdata,                --                .readdata
			m0_readdatavalid        => sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid,           --                .readdatavalid
			m0_read                 => sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent_m0_read,                    --                .read
			m0_waitrequest          => sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest,             --                .waitrequest
			m0_writedata            => sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent_m0_writedata,               --                .writedata
			m0_write                => sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent_m0_write,                   --                .write
			rp_endofpacket          => sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket,             --              rp.endofpacket
			rp_ready                => sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent_rp_ready,                   --                .ready
			rp_valid                => sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent_rp_valid,                   --                .valid
			rp_data                 => sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent_rp_data,                    --                .data
			rp_startofpacket        => sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket,           --                .startofpacket
			cp_ready                => cmd_xbar_demux_001_src3_ready,                                                                 --              cp.ready
			cp_valid                => cmd_xbar_demux_001_src3_valid,                                                                 --                .valid
			cp_data                 => cmd_xbar_demux_001_src3_data,                                                                  --                .data
			cp_startofpacket        => cmd_xbar_demux_001_src3_startofpacket,                                                         --                .startofpacket
			cp_endofpacket          => cmd_xbar_demux_001_src3_endofpacket,                                                           --                .endofpacket
			cp_channel              => cmd_xbar_demux_001_src3_channel,                                                               --                .channel
			rf_sink_ready           => sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready,         --         rf_sink.ready
			rf_sink_valid           => sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid,         --                .valid
			rf_sink_startofpacket   => sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket, --                .startofpacket
			rf_sink_endofpacket     => sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket,   --                .endofpacket
			rf_sink_data            => sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data,          --                .data
			rf_source_ready         => sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent_rf_source_ready,            --       rf_source.ready
			rf_source_valid         => sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent_rf_source_valid,            --                .valid
			rf_source_startofpacket => sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket,    --                .startofpacket
			rf_source_endofpacket   => sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket,      --                .endofpacket
			rf_source_data          => sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent_rf_source_data,             --                .data
			rdata_fifo_sink_ready   => sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready,       -- rdata_fifo_sink.ready
			rdata_fifo_sink_valid   => sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid,       --                .valid
			rdata_fifo_sink_data    => sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data,        --                .data
			rdata_fifo_src_ready    => sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready,       --  rdata_fifo_src.ready
			rdata_fifo_src_valid    => sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid,       --                .valid
			rdata_fifo_src_data     => sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data         --                .data
		);

	sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo : component Nios1_pio_LEDG_s1_translator_avalon_universal_slave_0_agent_rsp_fifo
		port map (
			clk               => clk_clk,                                                                                       --       clk.clk
			reset             => rst_controller_reset_out_reset,                                                                -- clk_reset.reset
			in_data           => sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent_rf_source_data,             --        in.data
			in_valid          => sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent_rf_source_valid,            --          .valid
			in_ready          => sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent_rf_source_ready,            --          .ready
			in_startofpacket  => sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket,    --          .startofpacket
			in_endofpacket    => sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket,      --          .endofpacket
			out_data          => sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data,          --       out.data
			out_valid         => sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid,         --          .valid
			out_ready         => sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready,         --          .ready
			out_startofpacket => sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket, --          .startofpacket
			out_endofpacket   => sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket    --          .endofpacket
		);

	pio_dataread_s1_translator_avalon_universal_slave_0_agent : component Nios1_pio_DataRead_s1_translator_avalon_universal_slave_0_agent
		port map (
			clk                     => clk_clk,                                                                              --             clk.clk
			reset                   => rst_controller_reset_out_reset,                                                       --       clk_reset.reset
			m0_address              => pio_dataread_s1_translator_avalon_universal_slave_0_agent_m0_address,                 --              m0.address
			m0_burstcount           => pio_dataread_s1_translator_avalon_universal_slave_0_agent_m0_burstcount,              --                .burstcount
			m0_byteenable           => pio_dataread_s1_translator_avalon_universal_slave_0_agent_m0_byteenable,              --                .byteenable
			m0_debugaccess          => pio_dataread_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess,             --                .debugaccess
			m0_lock                 => pio_dataread_s1_translator_avalon_universal_slave_0_agent_m0_lock,                    --                .lock
			m0_readdata             => pio_dataread_s1_translator_avalon_universal_slave_0_agent_m0_readdata,                --                .readdata
			m0_readdatavalid        => pio_dataread_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid,           --                .readdatavalid
			m0_read                 => pio_dataread_s1_translator_avalon_universal_slave_0_agent_m0_read,                    --                .read
			m0_waitrequest          => pio_dataread_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest,             --                .waitrequest
			m0_writedata            => pio_dataread_s1_translator_avalon_universal_slave_0_agent_m0_writedata,               --                .writedata
			m0_write                => pio_dataread_s1_translator_avalon_universal_slave_0_agent_m0_write,                   --                .write
			rp_endofpacket          => pio_dataread_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket,             --              rp.endofpacket
			rp_ready                => pio_dataread_s1_translator_avalon_universal_slave_0_agent_rp_ready,                   --                .ready
			rp_valid                => pio_dataread_s1_translator_avalon_universal_slave_0_agent_rp_valid,                   --                .valid
			rp_data                 => pio_dataread_s1_translator_avalon_universal_slave_0_agent_rp_data,                    --                .data
			rp_startofpacket        => pio_dataread_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket,           --                .startofpacket
			cp_ready                => cmd_xbar_demux_001_src13_ready,                                                       --              cp.ready
			cp_valid                => cmd_xbar_demux_001_src13_valid,                                                       --                .valid
			cp_data                 => cmd_xbar_demux_001_src13_data,                                                        --                .data
			cp_startofpacket        => cmd_xbar_demux_001_src13_startofpacket,                                               --                .startofpacket
			cp_endofpacket          => cmd_xbar_demux_001_src13_endofpacket,                                                 --                .endofpacket
			cp_channel              => cmd_xbar_demux_001_src13_channel,                                                     --                .channel
			rf_sink_ready           => pio_dataread_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready,         --         rf_sink.ready
			rf_sink_valid           => pio_dataread_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid,         --                .valid
			rf_sink_startofpacket   => pio_dataread_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket, --                .startofpacket
			rf_sink_endofpacket     => pio_dataread_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket,   --                .endofpacket
			rf_sink_data            => pio_dataread_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data,          --                .data
			rf_source_ready         => pio_dataread_s1_translator_avalon_universal_slave_0_agent_rf_source_ready,            --       rf_source.ready
			rf_source_valid         => pio_dataread_s1_translator_avalon_universal_slave_0_agent_rf_source_valid,            --                .valid
			rf_source_startofpacket => pio_dataread_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket,    --                .startofpacket
			rf_source_endofpacket   => pio_dataread_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket,      --                .endofpacket
			rf_source_data          => pio_dataread_s1_translator_avalon_universal_slave_0_agent_rf_source_data,             --                .data
			rdata_fifo_sink_ready   => pio_dataread_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready,       -- rdata_fifo_sink.ready
			rdata_fifo_sink_valid   => pio_dataread_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid,       --                .valid
			rdata_fifo_sink_data    => pio_dataread_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data,        --                .data
			rdata_fifo_src_ready    => pio_dataread_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready,       --  rdata_fifo_src.ready
			rdata_fifo_src_valid    => pio_dataread_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid,       --                .valid
			rdata_fifo_src_data     => pio_dataread_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data         --                .data
		);

	pio_dataread_s1_translator_avalon_universal_slave_0_agent_rsp_fifo : component Nios1_pio_LEDG_s1_translator_avalon_universal_slave_0_agent_rsp_fifo
		port map (
			clk               => clk_clk,                                                                              --       clk.clk
			reset             => rst_controller_reset_out_reset,                                                       -- clk_reset.reset
			in_data           => pio_dataread_s1_translator_avalon_universal_slave_0_agent_rf_source_data,             --        in.data
			in_valid          => pio_dataread_s1_translator_avalon_universal_slave_0_agent_rf_source_valid,            --          .valid
			in_ready          => pio_dataread_s1_translator_avalon_universal_slave_0_agent_rf_source_ready,            --          .ready
			in_startofpacket  => pio_dataread_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket,    --          .startofpacket
			in_endofpacket    => pio_dataread_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket,      --          .endofpacket
			out_data          => pio_dataread_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data,          --       out.data
			out_valid         => pio_dataread_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid,         --          .valid
			out_ready         => pio_dataread_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready,         --          .ready
			out_startofpacket => pio_dataread_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket, --          .startofpacket
			out_endofpacket   => pio_dataread_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket    --          .endofpacket
		);

	nios2_qsys_data_master_translator_avalon_universal_master_0_agent : component Nios1_nios2_qsys_data_master_translator_avalon_universal_master_0_agent
		port map (
			clk              => clk_clk,                                                                            --       clk.clk
			reset            => rst_controller_reset_out_reset,                                                     -- clk_reset.reset
			av_address       => nios2_qsys_data_master_translator_avalon_universal_master_0_address,                --        av.address
			av_write         => nios2_qsys_data_master_translator_avalon_universal_master_0_write,                  --          .write
			av_read          => nios2_qsys_data_master_translator_avalon_universal_master_0_read,                   --          .read
			av_writedata     => nios2_qsys_data_master_translator_avalon_universal_master_0_writedata,              --          .writedata
			av_readdata      => nios2_qsys_data_master_translator_avalon_universal_master_0_readdata,               --          .readdata
			av_waitrequest   => nios2_qsys_data_master_translator_avalon_universal_master_0_waitrequest,            --          .waitrequest
			av_readdatavalid => nios2_qsys_data_master_translator_avalon_universal_master_0_readdatavalid,          --          .readdatavalid
			av_byteenable    => nios2_qsys_data_master_translator_avalon_universal_master_0_byteenable,             --          .byteenable
			av_burstcount    => nios2_qsys_data_master_translator_avalon_universal_master_0_burstcount,             --          .burstcount
			av_debugaccess   => nios2_qsys_data_master_translator_avalon_universal_master_0_debugaccess,            --          .debugaccess
			av_lock          => nios2_qsys_data_master_translator_avalon_universal_master_0_lock,                   --          .lock
			cp_valid         => nios2_qsys_data_master_translator_avalon_universal_master_0_agent_cp_valid,         --        cp.valid
			cp_data          => nios2_qsys_data_master_translator_avalon_universal_master_0_agent_cp_data,          --          .data
			cp_startofpacket => nios2_qsys_data_master_translator_avalon_universal_master_0_agent_cp_startofpacket, --          .startofpacket
			cp_endofpacket   => nios2_qsys_data_master_translator_avalon_universal_master_0_agent_cp_endofpacket,   --          .endofpacket
			cp_ready         => nios2_qsys_data_master_translator_avalon_universal_master_0_agent_cp_ready,         --          .ready
			rp_valid         => limiter_001_rsp_src_valid,                                                          --        rp.valid
			rp_data          => limiter_001_rsp_src_data,                                                           --          .data
			rp_channel       => limiter_001_rsp_src_channel,                                                        --          .channel
			rp_startofpacket => limiter_001_rsp_src_startofpacket,                                                  --          .startofpacket
			rp_endofpacket   => limiter_001_rsp_src_endofpacket,                                                    --          .endofpacket
			rp_ready         => limiter_001_rsp_src_ready                                                           --          .ready
		);

	lcd_control_slave_translator_avalon_universal_slave_0_agent : component Nios1_lcd_control_slave_translator_avalon_universal_slave_0_agent
		port map (
			clk                     => clk_clk,                                                                                --             clk.clk
			reset                   => rst_controller_reset_out_reset,                                                         --       clk_reset.reset
			m0_address              => lcd_control_slave_translator_avalon_universal_slave_0_agent_m0_address,                 --              m0.address
			m0_burstcount           => lcd_control_slave_translator_avalon_universal_slave_0_agent_m0_burstcount,              --                .burstcount
			m0_byteenable           => lcd_control_slave_translator_avalon_universal_slave_0_agent_m0_byteenable,              --                .byteenable
			m0_debugaccess          => lcd_control_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess,             --                .debugaccess
			m0_lock                 => lcd_control_slave_translator_avalon_universal_slave_0_agent_m0_lock,                    --                .lock
			m0_readdata             => lcd_control_slave_translator_avalon_universal_slave_0_agent_m0_readdata,                --                .readdata
			m0_readdatavalid        => lcd_control_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid,           --                .readdatavalid
			m0_read                 => lcd_control_slave_translator_avalon_universal_slave_0_agent_m0_read,                    --                .read
			m0_waitrequest          => lcd_control_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest,             --                .waitrequest
			m0_writedata            => lcd_control_slave_translator_avalon_universal_slave_0_agent_m0_writedata,               --                .writedata
			m0_write                => lcd_control_slave_translator_avalon_universal_slave_0_agent_m0_write,                   --                .write
			rp_endofpacket          => lcd_control_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket,             --              rp.endofpacket
			rp_ready                => lcd_control_slave_translator_avalon_universal_slave_0_agent_rp_ready,                   --                .ready
			rp_valid                => lcd_control_slave_translator_avalon_universal_slave_0_agent_rp_valid,                   --                .valid
			rp_data                 => lcd_control_slave_translator_avalon_universal_slave_0_agent_rp_data,                    --                .data
			rp_startofpacket        => lcd_control_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket,           --                .startofpacket
			cp_ready                => cmd_xbar_demux_001_src8_ready,                                                          --              cp.ready
			cp_valid                => cmd_xbar_demux_001_src8_valid,                                                          --                .valid
			cp_data                 => cmd_xbar_demux_001_src8_data,                                                           --                .data
			cp_startofpacket        => cmd_xbar_demux_001_src8_startofpacket,                                                  --                .startofpacket
			cp_endofpacket          => cmd_xbar_demux_001_src8_endofpacket,                                                    --                .endofpacket
			cp_channel              => cmd_xbar_demux_001_src8_channel,                                                        --                .channel
			rf_sink_ready           => lcd_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready,         --         rf_sink.ready
			rf_sink_valid           => lcd_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid,         --                .valid
			rf_sink_startofpacket   => lcd_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket, --                .startofpacket
			rf_sink_endofpacket     => lcd_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket,   --                .endofpacket
			rf_sink_data            => lcd_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data,          --                .data
			rf_source_ready         => lcd_control_slave_translator_avalon_universal_slave_0_agent_rf_source_ready,            --       rf_source.ready
			rf_source_valid         => lcd_control_slave_translator_avalon_universal_slave_0_agent_rf_source_valid,            --                .valid
			rf_source_startofpacket => lcd_control_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket,    --                .startofpacket
			rf_source_endofpacket   => lcd_control_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket,      --                .endofpacket
			rf_source_data          => lcd_control_slave_translator_avalon_universal_slave_0_agent_rf_source_data,             --                .data
			rdata_fifo_sink_ready   => lcd_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready,       -- rdata_fifo_sink.ready
			rdata_fifo_sink_valid   => lcd_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid,       --                .valid
			rdata_fifo_sink_data    => lcd_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data,        --                .data
			rdata_fifo_src_ready    => lcd_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready,       --  rdata_fifo_src.ready
			rdata_fifo_src_valid    => lcd_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid,       --                .valid
			rdata_fifo_src_data     => lcd_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data         --                .data
		);

	lcd_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo : component Nios1_pio_LEDG_s1_translator_avalon_universal_slave_0_agent_rsp_fifo
		port map (
			clk               => clk_clk,                                                                                --       clk.clk
			reset             => rst_controller_reset_out_reset,                                                         -- clk_reset.reset
			in_data           => lcd_control_slave_translator_avalon_universal_slave_0_agent_rf_source_data,             --        in.data
			in_valid          => lcd_control_slave_translator_avalon_universal_slave_0_agent_rf_source_valid,            --          .valid
			in_ready          => lcd_control_slave_translator_avalon_universal_slave_0_agent_rf_source_ready,            --          .ready
			in_startofpacket  => lcd_control_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket,    --          .startofpacket
			in_endofpacket    => lcd_control_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket,      --          .endofpacket
			out_data          => lcd_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data,          --       out.data
			out_valid         => lcd_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid,         --          .valid
			out_ready         => lcd_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready,         --          .ready
			out_startofpacket => lcd_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket, --          .startofpacket
			out_endofpacket   => lcd_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket    --          .endofpacket
		);

	nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent : component Nios1_nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent
		port map (
			clk                     => clk_clk,                                                                                           --             clk.clk
			reset                   => rst_controller_reset_out_reset,                                                                    --       clk_reset.reset
			m0_address              => nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_address,                 --              m0.address
			m0_burstcount           => nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_burstcount,              --                .burstcount
			m0_byteenable           => nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_byteenable,              --                .byteenable
			m0_debugaccess          => nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_debugaccess,             --                .debugaccess
			m0_lock                 => nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_lock,                    --                .lock
			m0_readdata             => nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_readdata,                --                .readdata
			m0_readdatavalid        => nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_readdatavalid,           --                .readdatavalid
			m0_read                 => nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_read,                    --                .read
			m0_waitrequest          => nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_waitrequest,             --                .waitrequest
			m0_writedata            => nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_writedata,               --                .writedata
			m0_write                => nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_write,                   --                .write
			rp_endofpacket          => nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_endofpacket,             --              rp.endofpacket
			rp_ready                => nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_ready,                   --                .ready
			rp_valid                => nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_valid,                   --                .valid
			rp_data                 => nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_data,                    --                .data
			rp_startofpacket        => nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_startofpacket,           --                .startofpacket
			cp_ready                => cmd_xbar_mux_src_ready,                                                                            --              cp.ready
			cp_valid                => cmd_xbar_mux_src_valid,                                                                            --                .valid
			cp_data                 => cmd_xbar_mux_src_data,                                                                             --                .data
			cp_startofpacket        => cmd_xbar_mux_src_startofpacket,                                                                    --                .startofpacket
			cp_endofpacket          => cmd_xbar_mux_src_endofpacket,                                                                      --                .endofpacket
			cp_channel              => cmd_xbar_mux_src_channel,                                                                          --                .channel
			rf_sink_ready           => nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready,         --         rf_sink.ready
			rf_sink_valid           => nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid,         --                .valid
			rf_sink_startofpacket   => nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket, --                .startofpacket
			rf_sink_endofpacket     => nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket,   --                .endofpacket
			rf_sink_data            => nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data,          --                .data
			rf_source_ready         => nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_ready,            --       rf_source.ready
			rf_source_valid         => nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_valid,            --                .valid
			rf_source_startofpacket => nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_startofpacket,    --                .startofpacket
			rf_source_endofpacket   => nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_endofpacket,      --                .endofpacket
			rf_source_data          => nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_data,             --                .data
			rdata_fifo_sink_ready   => nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready,       -- rdata_fifo_sink.ready
			rdata_fifo_sink_valid   => nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid,       --                .valid
			rdata_fifo_sink_data    => nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data,        --                .data
			rdata_fifo_src_ready    => nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready,       --  rdata_fifo_src.ready
			rdata_fifo_src_valid    => nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid,       --                .valid
			rdata_fifo_src_data     => nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data         --                .data
		);

	nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo : component Nios1_pio_LEDG_s1_translator_avalon_universal_slave_0_agent_rsp_fifo
		port map (
			clk               => clk_clk,                                                                                           --       clk.clk
			reset             => rst_controller_reset_out_reset,                                                                    -- clk_reset.reset
			in_data           => nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_data,             --        in.data
			in_valid          => nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_valid,            --          .valid
			in_ready          => nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_ready,            --          .ready
			in_startofpacket  => nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_startofpacket,    --          .startofpacket
			in_endofpacket    => nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_endofpacket,      --          .endofpacket
			out_data          => nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data,          --       out.data
			out_valid         => nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid,         --          .valid
			out_ready         => nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready,         --          .ready
			out_startofpacket => nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket, --          .startofpacket
			out_endofpacket   => nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket    --          .endofpacket
		);

	nios2_qsys_instruction_master_translator_avalon_universal_master_0_agent : component Nios1_nios2_qsys_instruction_master_translator_avalon_universal_master_0_agent
		port map (
			clk              => clk_clk,                                                                                   --       clk.clk
			reset            => rst_controller_reset_out_reset,                                                            -- clk_reset.reset
			av_address       => nios2_qsys_instruction_master_translator_avalon_universal_master_0_address,                --        av.address
			av_write         => nios2_qsys_instruction_master_translator_avalon_universal_master_0_write,                  --          .write
			av_read          => nios2_qsys_instruction_master_translator_avalon_universal_master_0_read,                   --          .read
			av_writedata     => nios2_qsys_instruction_master_translator_avalon_universal_master_0_writedata,              --          .writedata
			av_readdata      => nios2_qsys_instruction_master_translator_avalon_universal_master_0_readdata,               --          .readdata
			av_waitrequest   => nios2_qsys_instruction_master_translator_avalon_universal_master_0_waitrequest,            --          .waitrequest
			av_readdatavalid => nios2_qsys_instruction_master_translator_avalon_universal_master_0_readdatavalid,          --          .readdatavalid
			av_byteenable    => nios2_qsys_instruction_master_translator_avalon_universal_master_0_byteenable,             --          .byteenable
			av_burstcount    => nios2_qsys_instruction_master_translator_avalon_universal_master_0_burstcount,             --          .burstcount
			av_debugaccess   => nios2_qsys_instruction_master_translator_avalon_universal_master_0_debugaccess,            --          .debugaccess
			av_lock          => nios2_qsys_instruction_master_translator_avalon_universal_master_0_lock,                   --          .lock
			cp_valid         => nios2_qsys_instruction_master_translator_avalon_universal_master_0_agent_cp_valid,         --        cp.valid
			cp_data          => nios2_qsys_instruction_master_translator_avalon_universal_master_0_agent_cp_data,          --          .data
			cp_startofpacket => nios2_qsys_instruction_master_translator_avalon_universal_master_0_agent_cp_startofpacket, --          .startofpacket
			cp_endofpacket   => nios2_qsys_instruction_master_translator_avalon_universal_master_0_agent_cp_endofpacket,   --          .endofpacket
			cp_ready         => nios2_qsys_instruction_master_translator_avalon_universal_master_0_agent_cp_ready,         --          .ready
			rp_valid         => limiter_rsp_src_valid,                                                                     --        rp.valid
			rp_data          => limiter_rsp_src_data,                                                                      --          .data
			rp_channel       => limiter_rsp_src_channel,                                                                   --          .channel
			rp_startofpacket => limiter_rsp_src_startofpacket,                                                             --          .startofpacket
			rp_endofpacket   => limiter_rsp_src_endofpacket,                                                               --          .endofpacket
			rp_ready         => limiter_rsp_src_ready                                                                      --          .ready
		);

	pio_sw_s1_translator_avalon_universal_slave_0_agent : component Nios1_pio_SW_s1_translator_avalon_universal_slave_0_agent
		port map (
			clk                     => clk_clk,                                                                        --             clk.clk
			reset                   => rst_controller_reset_out_reset,                                                 --       clk_reset.reset
			m0_address              => pio_sw_s1_translator_avalon_universal_slave_0_agent_m0_address,                 --              m0.address
			m0_burstcount           => pio_sw_s1_translator_avalon_universal_slave_0_agent_m0_burstcount,              --                .burstcount
			m0_byteenable           => pio_sw_s1_translator_avalon_universal_slave_0_agent_m0_byteenable,              --                .byteenable
			m0_debugaccess          => pio_sw_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess,             --                .debugaccess
			m0_lock                 => pio_sw_s1_translator_avalon_universal_slave_0_agent_m0_lock,                    --                .lock
			m0_readdata             => pio_sw_s1_translator_avalon_universal_slave_0_agent_m0_readdata,                --                .readdata
			m0_readdatavalid        => pio_sw_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid,           --                .readdatavalid
			m0_read                 => pio_sw_s1_translator_avalon_universal_slave_0_agent_m0_read,                    --                .read
			m0_waitrequest          => pio_sw_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest,             --                .waitrequest
			m0_writedata            => pio_sw_s1_translator_avalon_universal_slave_0_agent_m0_writedata,               --                .writedata
			m0_write                => pio_sw_s1_translator_avalon_universal_slave_0_agent_m0_write,                   --                .write
			rp_endofpacket          => pio_sw_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket,             --              rp.endofpacket
			rp_ready                => pio_sw_s1_translator_avalon_universal_slave_0_agent_rp_ready,                   --                .ready
			rp_valid                => pio_sw_s1_translator_avalon_universal_slave_0_agent_rp_valid,                   --                .valid
			rp_data                 => pio_sw_s1_translator_avalon_universal_slave_0_agent_rp_data,                    --                .data
			rp_startofpacket        => pio_sw_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket,           --                .startofpacket
			cp_ready                => cmd_xbar_demux_001_src6_ready,                                                  --              cp.ready
			cp_valid                => cmd_xbar_demux_001_src6_valid,                                                  --                .valid
			cp_data                 => cmd_xbar_demux_001_src6_data,                                                   --                .data
			cp_startofpacket        => cmd_xbar_demux_001_src6_startofpacket,                                          --                .startofpacket
			cp_endofpacket          => cmd_xbar_demux_001_src6_endofpacket,                                            --                .endofpacket
			cp_channel              => cmd_xbar_demux_001_src6_channel,                                                --                .channel
			rf_sink_ready           => pio_sw_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready,         --         rf_sink.ready
			rf_sink_valid           => pio_sw_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid,         --                .valid
			rf_sink_startofpacket   => pio_sw_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket, --                .startofpacket
			rf_sink_endofpacket     => pio_sw_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket,   --                .endofpacket
			rf_sink_data            => pio_sw_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data,          --                .data
			rf_source_ready         => pio_sw_s1_translator_avalon_universal_slave_0_agent_rf_source_ready,            --       rf_source.ready
			rf_source_valid         => pio_sw_s1_translator_avalon_universal_slave_0_agent_rf_source_valid,            --                .valid
			rf_source_startofpacket => pio_sw_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket,    --                .startofpacket
			rf_source_endofpacket   => pio_sw_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket,      --                .endofpacket
			rf_source_data          => pio_sw_s1_translator_avalon_universal_slave_0_agent_rf_source_data,             --                .data
			rdata_fifo_sink_ready   => pio_sw_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready,       -- rdata_fifo_sink.ready
			rdata_fifo_sink_valid   => pio_sw_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid,       --                .valid
			rdata_fifo_sink_data    => pio_sw_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data,        --                .data
			rdata_fifo_src_ready    => pio_sw_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready,       --  rdata_fifo_src.ready
			rdata_fifo_src_valid    => pio_sw_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid,       --                .valid
			rdata_fifo_src_data     => pio_sw_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data         --                .data
		);

	pio_sw_s1_translator_avalon_universal_slave_0_agent_rsp_fifo : component Nios1_pio_LEDG_s1_translator_avalon_universal_slave_0_agent_rsp_fifo
		port map (
			clk               => clk_clk,                                                                        --       clk.clk
			reset             => rst_controller_reset_out_reset,                                                 -- clk_reset.reset
			in_data           => pio_sw_s1_translator_avalon_universal_slave_0_agent_rf_source_data,             --        in.data
			in_valid          => pio_sw_s1_translator_avalon_universal_slave_0_agent_rf_source_valid,            --          .valid
			in_ready          => pio_sw_s1_translator_avalon_universal_slave_0_agent_rf_source_ready,            --          .ready
			in_startofpacket  => pio_sw_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket,    --          .startofpacket
			in_endofpacket    => pio_sw_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket,      --          .endofpacket
			out_data          => pio_sw_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data,          --       out.data
			out_valid         => pio_sw_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid,         --          .valid
			out_ready         => pio_sw_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready,         --          .ready
			out_startofpacket => pio_sw_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket, --          .startofpacket
			out_endofpacket   => pio_sw_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket    --          .endofpacket
		);

	jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent : component Nios1_jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent
		port map (
			clk                     => clk_clk,                                                                                          --             clk.clk
			reset                   => rst_controller_reset_out_reset,                                                                   --       clk_reset.reset
			m0_address              => jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_address,                 --              m0.address
			m0_burstcount           => jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_burstcount,              --                .burstcount
			m0_byteenable           => jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_byteenable,              --                .byteenable
			m0_debugaccess          => jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess,             --                .debugaccess
			m0_lock                 => jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_lock,                    --                .lock
			m0_readdata             => jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_readdata,                --                .readdata
			m0_readdatavalid        => jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid,           --                .readdatavalid
			m0_read                 => jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_read,                    --                .read
			m0_waitrequest          => jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest,             --                .waitrequest
			m0_writedata            => jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_writedata,               --                .writedata
			m0_write                => jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_write,                   --                .write
			rp_endofpacket          => jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket,             --              rp.endofpacket
			rp_ready                => jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_ready,                   --                .ready
			rp_valid                => jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_valid,                   --                .valid
			rp_data                 => jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_data,                    --                .data
			rp_startofpacket        => jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket,           --                .startofpacket
			cp_ready                => cmd_xbar_demux_001_src2_ready,                                                                    --              cp.ready
			cp_valid                => cmd_xbar_demux_001_src2_valid,                                                                    --                .valid
			cp_data                 => cmd_xbar_demux_001_src2_data,                                                                     --                .data
			cp_startofpacket        => cmd_xbar_demux_001_src2_startofpacket,                                                            --                .startofpacket
			cp_endofpacket          => cmd_xbar_demux_001_src2_endofpacket,                                                              --                .endofpacket
			cp_channel              => cmd_xbar_demux_001_src2_channel,                                                                  --                .channel
			rf_sink_ready           => jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready,         --         rf_sink.ready
			rf_sink_valid           => jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid,         --                .valid
			rf_sink_startofpacket   => jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket, --                .startofpacket
			rf_sink_endofpacket     => jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket,   --                .endofpacket
			rf_sink_data            => jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data,          --                .data
			rf_source_ready         => jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_ready,            --       rf_source.ready
			rf_source_valid         => jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_valid,            --                .valid
			rf_source_startofpacket => jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket,    --                .startofpacket
			rf_source_endofpacket   => jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket,      --                .endofpacket
			rf_source_data          => jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_data,             --                .data
			rdata_fifo_sink_ready   => jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready,       -- rdata_fifo_sink.ready
			rdata_fifo_sink_valid   => jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid,       --                .valid
			rdata_fifo_sink_data    => jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data,        --                .data
			rdata_fifo_src_ready    => jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready,       --  rdata_fifo_src.ready
			rdata_fifo_src_valid    => jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid,       --                .valid
			rdata_fifo_src_data     => jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data         --                .data
		);

	jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo : component Nios1_pio_LEDG_s1_translator_avalon_universal_slave_0_agent_rsp_fifo
		port map (
			clk               => clk_clk,                                                                                          --       clk.clk
			reset             => rst_controller_reset_out_reset,                                                                   -- clk_reset.reset
			in_data           => jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_data,             --        in.data
			in_valid          => jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_valid,            --          .valid
			in_ready          => jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_ready,            --          .ready
			in_startofpacket  => jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket,    --          .startofpacket
			in_endofpacket    => jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket,      --          .endofpacket
			out_data          => jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data,          --       out.data
			out_valid         => jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid,         --          .valid
			out_ready         => jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready,         --          .ready
			out_startofpacket => jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket, --          .startofpacket
			out_endofpacket   => jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket    --          .endofpacket
		);

	pio_button_s1_translator_avalon_universal_slave_0_agent : component Nios1_pio_Button_s1_translator_avalon_universal_slave_0_agent
		port map (
			clk                     => clk_clk,                                                                            --             clk.clk
			reset                   => rst_controller_reset_out_reset,                                                     --       clk_reset.reset
			m0_address              => pio_button_s1_translator_avalon_universal_slave_0_agent_m0_address,                 --              m0.address
			m0_burstcount           => pio_button_s1_translator_avalon_universal_slave_0_agent_m0_burstcount,              --                .burstcount
			m0_byteenable           => pio_button_s1_translator_avalon_universal_slave_0_agent_m0_byteenable,              --                .byteenable
			m0_debugaccess          => pio_button_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess,             --                .debugaccess
			m0_lock                 => pio_button_s1_translator_avalon_universal_slave_0_agent_m0_lock,                    --                .lock
			m0_readdata             => pio_button_s1_translator_avalon_universal_slave_0_agent_m0_readdata,                --                .readdata
			m0_readdatavalid        => pio_button_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid,           --                .readdatavalid
			m0_read                 => pio_button_s1_translator_avalon_universal_slave_0_agent_m0_read,                    --                .read
			m0_waitrequest          => pio_button_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest,             --                .waitrequest
			m0_writedata            => pio_button_s1_translator_avalon_universal_slave_0_agent_m0_writedata,               --                .writedata
			m0_write                => pio_button_s1_translator_avalon_universal_slave_0_agent_m0_write,                   --                .write
			rp_endofpacket          => pio_button_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket,             --              rp.endofpacket
			rp_ready                => pio_button_s1_translator_avalon_universal_slave_0_agent_rp_ready,                   --                .ready
			rp_valid                => pio_button_s1_translator_avalon_universal_slave_0_agent_rp_valid,                   --                .valid
			rp_data                 => pio_button_s1_translator_avalon_universal_slave_0_agent_rp_data,                    --                .data
			rp_startofpacket        => pio_button_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket,           --                .startofpacket
			cp_ready                => cmd_xbar_demux_001_src7_ready,                                                      --              cp.ready
			cp_valid                => cmd_xbar_demux_001_src7_valid,                                                      --                .valid
			cp_data                 => cmd_xbar_demux_001_src7_data,                                                       --                .data
			cp_startofpacket        => cmd_xbar_demux_001_src7_startofpacket,                                              --                .startofpacket
			cp_endofpacket          => cmd_xbar_demux_001_src7_endofpacket,                                                --                .endofpacket
			cp_channel              => cmd_xbar_demux_001_src7_channel,                                                    --                .channel
			rf_sink_ready           => pio_button_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready,         --         rf_sink.ready
			rf_sink_valid           => pio_button_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid,         --                .valid
			rf_sink_startofpacket   => pio_button_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket, --                .startofpacket
			rf_sink_endofpacket     => pio_button_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket,   --                .endofpacket
			rf_sink_data            => pio_button_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data,          --                .data
			rf_source_ready         => pio_button_s1_translator_avalon_universal_slave_0_agent_rf_source_ready,            --       rf_source.ready
			rf_source_valid         => pio_button_s1_translator_avalon_universal_slave_0_agent_rf_source_valid,            --                .valid
			rf_source_startofpacket => pio_button_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket,    --                .startofpacket
			rf_source_endofpacket   => pio_button_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket,      --                .endofpacket
			rf_source_data          => pio_button_s1_translator_avalon_universal_slave_0_agent_rf_source_data,             --                .data
			rdata_fifo_sink_ready   => pio_button_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready,       -- rdata_fifo_sink.ready
			rdata_fifo_sink_valid   => pio_button_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid,       --                .valid
			rdata_fifo_sink_data    => pio_button_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data,        --                .data
			rdata_fifo_src_ready    => pio_button_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready,       --  rdata_fifo_src.ready
			rdata_fifo_src_valid    => pio_button_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid,       --                .valid
			rdata_fifo_src_data     => pio_button_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data         --                .data
		);

	pio_button_s1_translator_avalon_universal_slave_0_agent_rsp_fifo : component Nios1_pio_LEDG_s1_translator_avalon_universal_slave_0_agent_rsp_fifo
		port map (
			clk               => clk_clk,                                                                            --       clk.clk
			reset             => rst_controller_reset_out_reset,                                                     -- clk_reset.reset
			in_data           => pio_button_s1_translator_avalon_universal_slave_0_agent_rf_source_data,             --        in.data
			in_valid          => pio_button_s1_translator_avalon_universal_slave_0_agent_rf_source_valid,            --          .valid
			in_ready          => pio_button_s1_translator_avalon_universal_slave_0_agent_rf_source_ready,            --          .ready
			in_startofpacket  => pio_button_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket,    --          .startofpacket
			in_endofpacket    => pio_button_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket,      --          .endofpacket
			out_data          => pio_button_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data,          --       out.data
			out_valid         => pio_button_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid,         --          .valid
			out_ready         => pio_button_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready,         --          .ready
			out_startofpacket => pio_button_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket, --          .startofpacket
			out_endofpacket   => pio_button_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket    --          .endofpacket
		);

	pio_data_s1_translator_avalon_universal_slave_0_agent : component Nios1_pio_Data_s1_translator_avalon_universal_slave_0_agent
		port map (
			clk                     => clk_clk,                                                                          --             clk.clk
			reset                   => rst_controller_reset_out_reset,                                                   --       clk_reset.reset
			m0_address              => pio_data_s1_translator_avalon_universal_slave_0_agent_m0_address,                 --              m0.address
			m0_burstcount           => pio_data_s1_translator_avalon_universal_slave_0_agent_m0_burstcount,              --                .burstcount
			m0_byteenable           => pio_data_s1_translator_avalon_universal_slave_0_agent_m0_byteenable,              --                .byteenable
			m0_debugaccess          => pio_data_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess,             --                .debugaccess
			m0_lock                 => pio_data_s1_translator_avalon_universal_slave_0_agent_m0_lock,                    --                .lock
			m0_readdata             => pio_data_s1_translator_avalon_universal_slave_0_agent_m0_readdata,                --                .readdata
			m0_readdatavalid        => pio_data_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid,           --                .readdatavalid
			m0_read                 => pio_data_s1_translator_avalon_universal_slave_0_agent_m0_read,                    --                .read
			m0_waitrequest          => pio_data_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest,             --                .waitrequest
			m0_writedata            => pio_data_s1_translator_avalon_universal_slave_0_agent_m0_writedata,               --                .writedata
			m0_write                => pio_data_s1_translator_avalon_universal_slave_0_agent_m0_write,                   --                .write
			rp_endofpacket          => pio_data_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket,             --              rp.endofpacket
			rp_ready                => pio_data_s1_translator_avalon_universal_slave_0_agent_rp_ready,                   --                .ready
			rp_valid                => pio_data_s1_translator_avalon_universal_slave_0_agent_rp_valid,                   --                .valid
			rp_data                 => pio_data_s1_translator_avalon_universal_slave_0_agent_rp_data,                    --                .data
			rp_startofpacket        => pio_data_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket,           --                .startofpacket
			cp_ready                => cmd_xbar_demux_001_src11_ready,                                                   --              cp.ready
			cp_valid                => cmd_xbar_demux_001_src11_valid,                                                   --                .valid
			cp_data                 => cmd_xbar_demux_001_src11_data,                                                    --                .data
			cp_startofpacket        => cmd_xbar_demux_001_src11_startofpacket,                                           --                .startofpacket
			cp_endofpacket          => cmd_xbar_demux_001_src11_endofpacket,                                             --                .endofpacket
			cp_channel              => cmd_xbar_demux_001_src11_channel,                                                 --                .channel
			rf_sink_ready           => pio_data_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready,         --         rf_sink.ready
			rf_sink_valid           => pio_data_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid,         --                .valid
			rf_sink_startofpacket   => pio_data_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket, --                .startofpacket
			rf_sink_endofpacket     => pio_data_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket,   --                .endofpacket
			rf_sink_data            => pio_data_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data,          --                .data
			rf_source_ready         => pio_data_s1_translator_avalon_universal_slave_0_agent_rf_source_ready,            --       rf_source.ready
			rf_source_valid         => pio_data_s1_translator_avalon_universal_slave_0_agent_rf_source_valid,            --                .valid
			rf_source_startofpacket => pio_data_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket,    --                .startofpacket
			rf_source_endofpacket   => pio_data_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket,      --                .endofpacket
			rf_source_data          => pio_data_s1_translator_avalon_universal_slave_0_agent_rf_source_data,             --                .data
			rdata_fifo_sink_ready   => pio_data_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready,       -- rdata_fifo_sink.ready
			rdata_fifo_sink_valid   => pio_data_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid,       --                .valid
			rdata_fifo_sink_data    => pio_data_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data,        --                .data
			rdata_fifo_src_ready    => pio_data_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready,       --  rdata_fifo_src.ready
			rdata_fifo_src_valid    => pio_data_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid,       --                .valid
			rdata_fifo_src_data     => pio_data_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data         --                .data
		);

	pio_data_s1_translator_avalon_universal_slave_0_agent_rsp_fifo : component Nios1_pio_LEDG_s1_translator_avalon_universal_slave_0_agent_rsp_fifo
		port map (
			clk               => clk_clk,                                                                          --       clk.clk
			reset             => rst_controller_reset_out_reset,                                                   -- clk_reset.reset
			in_data           => pio_data_s1_translator_avalon_universal_slave_0_agent_rf_source_data,             --        in.data
			in_valid          => pio_data_s1_translator_avalon_universal_slave_0_agent_rf_source_valid,            --          .valid
			in_ready          => pio_data_s1_translator_avalon_universal_slave_0_agent_rf_source_ready,            --          .ready
			in_startofpacket  => pio_data_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket,    --          .startofpacket
			in_endofpacket    => pio_data_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket,      --          .endofpacket
			out_data          => pio_data_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data,          --       out.data
			out_valid         => pio_data_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid,         --          .valid
			out_ready         => pio_data_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready,         --          .ready
			out_startofpacket => pio_data_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket, --          .startofpacket
			out_endofpacket   => pio_data_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket    --          .endofpacket
		);

	uart_s1_translator_avalon_universal_slave_0_agent : component Nios1_uart_s1_translator_avalon_universal_slave_0_agent
		port map (
			clk                     => clk_clk,                                                                      --             clk.clk
			reset                   => rst_controller_reset_out_reset,                                               --       clk_reset.reset
			m0_address              => uart_s1_translator_avalon_universal_slave_0_agent_m0_address,                 --              m0.address
			m0_burstcount           => uart_s1_translator_avalon_universal_slave_0_agent_m0_burstcount,              --                .burstcount
			m0_byteenable           => uart_s1_translator_avalon_universal_slave_0_agent_m0_byteenable,              --                .byteenable
			m0_debugaccess          => uart_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess,             --                .debugaccess
			m0_lock                 => uart_s1_translator_avalon_universal_slave_0_agent_m0_lock,                    --                .lock
			m0_readdata             => uart_s1_translator_avalon_universal_slave_0_agent_m0_readdata,                --                .readdata
			m0_readdatavalid        => uart_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid,           --                .readdatavalid
			m0_read                 => uart_s1_translator_avalon_universal_slave_0_agent_m0_read,                    --                .read
			m0_waitrequest          => uart_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest,             --                .waitrequest
			m0_writedata            => uart_s1_translator_avalon_universal_slave_0_agent_m0_writedata,               --                .writedata
			m0_write                => uart_s1_translator_avalon_universal_slave_0_agent_m0_write,                   --                .write
			rp_endofpacket          => uart_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket,             --              rp.endofpacket
			rp_ready                => uart_s1_translator_avalon_universal_slave_0_agent_rp_ready,                   --                .ready
			rp_valid                => uart_s1_translator_avalon_universal_slave_0_agent_rp_valid,                   --                .valid
			rp_data                 => uart_s1_translator_avalon_universal_slave_0_agent_rp_data,                    --                .data
			rp_startofpacket        => uart_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket,           --                .startofpacket
			cp_ready                => cmd_xbar_demux_001_src9_ready,                                                --              cp.ready
			cp_valid                => cmd_xbar_demux_001_src9_valid,                                                --                .valid
			cp_data                 => cmd_xbar_demux_001_src9_data,                                                 --                .data
			cp_startofpacket        => cmd_xbar_demux_001_src9_startofpacket,                                        --                .startofpacket
			cp_endofpacket          => cmd_xbar_demux_001_src9_endofpacket,                                          --                .endofpacket
			cp_channel              => cmd_xbar_demux_001_src9_channel,                                              --                .channel
			rf_sink_ready           => uart_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready,         --         rf_sink.ready
			rf_sink_valid           => uart_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid,         --                .valid
			rf_sink_startofpacket   => uart_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket, --                .startofpacket
			rf_sink_endofpacket     => uart_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket,   --                .endofpacket
			rf_sink_data            => uart_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data,          --                .data
			rf_source_ready         => uart_s1_translator_avalon_universal_slave_0_agent_rf_source_ready,            --       rf_source.ready
			rf_source_valid         => uart_s1_translator_avalon_universal_slave_0_agent_rf_source_valid,            --                .valid
			rf_source_startofpacket => uart_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket,    --                .startofpacket
			rf_source_endofpacket   => uart_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket,      --                .endofpacket
			rf_source_data          => uart_s1_translator_avalon_universal_slave_0_agent_rf_source_data,             --                .data
			rdata_fifo_sink_ready   => uart_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready,       -- rdata_fifo_sink.ready
			rdata_fifo_sink_valid   => uart_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid,       --                .valid
			rdata_fifo_sink_data    => uart_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data,        --                .data
			rdata_fifo_src_ready    => uart_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready,       --  rdata_fifo_src.ready
			rdata_fifo_src_valid    => uart_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid,       --                .valid
			rdata_fifo_src_data     => uart_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data         --                .data
		);

	uart_s1_translator_avalon_universal_slave_0_agent_rsp_fifo : component Nios1_pio_LEDG_s1_translator_avalon_universal_slave_0_agent_rsp_fifo
		port map (
			clk               => clk_clk,                                                                      --       clk.clk
			reset             => rst_controller_reset_out_reset,                                               -- clk_reset.reset
			in_data           => uart_s1_translator_avalon_universal_slave_0_agent_rf_source_data,             --        in.data
			in_valid          => uart_s1_translator_avalon_universal_slave_0_agent_rf_source_valid,            --          .valid
			in_ready          => uart_s1_translator_avalon_universal_slave_0_agent_rf_source_ready,            --          .ready
			in_startofpacket  => uart_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket,    --          .startofpacket
			in_endofpacket    => uart_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket,      --          .endofpacket
			out_data          => uart_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data,          --       out.data
			out_valid         => uart_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid,         --          .valid
			out_ready         => uart_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready,         --          .ready
			out_startofpacket => uart_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket, --          .startofpacket
			out_endofpacket   => uart_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket    --          .endofpacket
		);

	onchip_memory_s1_translator_avalon_universal_slave_0_agent : component Nios1_onchip_memory_s1_translator_avalon_universal_slave_0_agent
		port map (
			clk                     => clk_clk,                                                                               --             clk.clk
			reset                   => rst_controller_reset_out_reset,                                                        --       clk_reset.reset
			m0_address              => onchip_memory_s1_translator_avalon_universal_slave_0_agent_m0_address,                 --              m0.address
			m0_burstcount           => onchip_memory_s1_translator_avalon_universal_slave_0_agent_m0_burstcount,              --                .burstcount
			m0_byteenable           => onchip_memory_s1_translator_avalon_universal_slave_0_agent_m0_byteenable,              --                .byteenable
			m0_debugaccess          => onchip_memory_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess,             --                .debugaccess
			m0_lock                 => onchip_memory_s1_translator_avalon_universal_slave_0_agent_m0_lock,                    --                .lock
			m0_readdata             => onchip_memory_s1_translator_avalon_universal_slave_0_agent_m0_readdata,                --                .readdata
			m0_readdatavalid        => onchip_memory_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid,           --                .readdatavalid
			m0_read                 => onchip_memory_s1_translator_avalon_universal_slave_0_agent_m0_read,                    --                .read
			m0_waitrequest          => onchip_memory_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest,             --                .waitrequest
			m0_writedata            => onchip_memory_s1_translator_avalon_universal_slave_0_agent_m0_writedata,               --                .writedata
			m0_write                => onchip_memory_s1_translator_avalon_universal_slave_0_agent_m0_write,                   --                .write
			rp_endofpacket          => onchip_memory_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket,             --              rp.endofpacket
			rp_ready                => onchip_memory_s1_translator_avalon_universal_slave_0_agent_rp_ready,                   --                .ready
			rp_valid                => onchip_memory_s1_translator_avalon_universal_slave_0_agent_rp_valid,                   --                .valid
			rp_data                 => onchip_memory_s1_translator_avalon_universal_slave_0_agent_rp_data,                    --                .data
			rp_startofpacket        => onchip_memory_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket,           --                .startofpacket
			cp_ready                => cmd_xbar_mux_001_src_ready,                                                            --              cp.ready
			cp_valid                => cmd_xbar_mux_001_src_valid,                                                            --                .valid
			cp_data                 => cmd_xbar_mux_001_src_data,                                                             --                .data
			cp_startofpacket        => cmd_xbar_mux_001_src_startofpacket,                                                    --                .startofpacket
			cp_endofpacket          => cmd_xbar_mux_001_src_endofpacket,                                                      --                .endofpacket
			cp_channel              => cmd_xbar_mux_001_src_channel,                                                          --                .channel
			rf_sink_ready           => onchip_memory_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready,         --         rf_sink.ready
			rf_sink_valid           => onchip_memory_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid,         --                .valid
			rf_sink_startofpacket   => onchip_memory_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket, --                .startofpacket
			rf_sink_endofpacket     => onchip_memory_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket,   --                .endofpacket
			rf_sink_data            => onchip_memory_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data,          --                .data
			rf_source_ready         => onchip_memory_s1_translator_avalon_universal_slave_0_agent_rf_source_ready,            --       rf_source.ready
			rf_source_valid         => onchip_memory_s1_translator_avalon_universal_slave_0_agent_rf_source_valid,            --                .valid
			rf_source_startofpacket => onchip_memory_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket,    --                .startofpacket
			rf_source_endofpacket   => onchip_memory_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket,      --                .endofpacket
			rf_source_data          => onchip_memory_s1_translator_avalon_universal_slave_0_agent_rf_source_data,             --                .data
			rdata_fifo_sink_ready   => onchip_memory_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready,       -- rdata_fifo_sink.ready
			rdata_fifo_sink_valid   => onchip_memory_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid,       --                .valid
			rdata_fifo_sink_data    => onchip_memory_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data,        --                .data
			rdata_fifo_src_ready    => onchip_memory_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready,       --  rdata_fifo_src.ready
			rdata_fifo_src_valid    => onchip_memory_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid,       --                .valid
			rdata_fifo_src_data     => onchip_memory_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data         --                .data
		);

	onchip_memory_s1_translator_avalon_universal_slave_0_agent_rsp_fifo : component Nios1_pio_LEDG_s1_translator_avalon_universal_slave_0_agent_rsp_fifo
		port map (
			clk               => clk_clk,                                                                               --       clk.clk
			reset             => rst_controller_reset_out_reset,                                                        -- clk_reset.reset
			in_data           => onchip_memory_s1_translator_avalon_universal_slave_0_agent_rf_source_data,             --        in.data
			in_valid          => onchip_memory_s1_translator_avalon_universal_slave_0_agent_rf_source_valid,            --          .valid
			in_ready          => onchip_memory_s1_translator_avalon_universal_slave_0_agent_rf_source_ready,            --          .ready
			in_startofpacket  => onchip_memory_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket,    --          .startofpacket
			in_endofpacket    => onchip_memory_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket,      --          .endofpacket
			out_data          => onchip_memory_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data,          --       out.data
			out_valid         => onchip_memory_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid,         --          .valid
			out_ready         => onchip_memory_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready,         --          .ready
			out_startofpacket => onchip_memory_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket, --          .startofpacket
			out_endofpacket   => onchip_memory_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket    --          .endofpacket
		);

	timer_0_s1_translator_avalon_universal_slave_0_agent : component Nios1_timer_0_s1_translator_avalon_universal_slave_0_agent
		port map (
			clk                     => clk_clk,                                                                         --             clk.clk
			reset                   => rst_controller_reset_out_reset,                                                  --       clk_reset.reset
			m0_address              => timer_0_s1_translator_avalon_universal_slave_0_agent_m0_address,                 --              m0.address
			m0_burstcount           => timer_0_s1_translator_avalon_universal_slave_0_agent_m0_burstcount,              --                .burstcount
			m0_byteenable           => timer_0_s1_translator_avalon_universal_slave_0_agent_m0_byteenable,              --                .byteenable
			m0_debugaccess          => timer_0_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess,             --                .debugaccess
			m0_lock                 => timer_0_s1_translator_avalon_universal_slave_0_agent_m0_lock,                    --                .lock
			m0_readdata             => timer_0_s1_translator_avalon_universal_slave_0_agent_m0_readdata,                --                .readdata
			m0_readdatavalid        => timer_0_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid,           --                .readdatavalid
			m0_read                 => timer_0_s1_translator_avalon_universal_slave_0_agent_m0_read,                    --                .read
			m0_waitrequest          => timer_0_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest,             --                .waitrequest
			m0_writedata            => timer_0_s1_translator_avalon_universal_slave_0_agent_m0_writedata,               --                .writedata
			m0_write                => timer_0_s1_translator_avalon_universal_slave_0_agent_m0_write,                   --                .write
			rp_endofpacket          => timer_0_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket,             --              rp.endofpacket
			rp_ready                => timer_0_s1_translator_avalon_universal_slave_0_agent_rp_ready,                   --                .ready
			rp_valid                => timer_0_s1_translator_avalon_universal_slave_0_agent_rp_valid,                   --                .valid
			rp_data                 => timer_0_s1_translator_avalon_universal_slave_0_agent_rp_data,                    --                .data
			rp_startofpacket        => timer_0_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket,           --                .startofpacket
			cp_ready                => cmd_xbar_demux_001_src10_ready,                                                  --              cp.ready
			cp_valid                => cmd_xbar_demux_001_src10_valid,                                                  --                .valid
			cp_data                 => cmd_xbar_demux_001_src10_data,                                                   --                .data
			cp_startofpacket        => cmd_xbar_demux_001_src10_startofpacket,                                          --                .startofpacket
			cp_endofpacket          => cmd_xbar_demux_001_src10_endofpacket,                                            --                .endofpacket
			cp_channel              => cmd_xbar_demux_001_src10_channel,                                                --                .channel
			rf_sink_ready           => timer_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready,         --         rf_sink.ready
			rf_sink_valid           => timer_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid,         --                .valid
			rf_sink_startofpacket   => timer_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket, --                .startofpacket
			rf_sink_endofpacket     => timer_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket,   --                .endofpacket
			rf_sink_data            => timer_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data,          --                .data
			rf_source_ready         => timer_0_s1_translator_avalon_universal_slave_0_agent_rf_source_ready,            --       rf_source.ready
			rf_source_valid         => timer_0_s1_translator_avalon_universal_slave_0_agent_rf_source_valid,            --                .valid
			rf_source_startofpacket => timer_0_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket,    --                .startofpacket
			rf_source_endofpacket   => timer_0_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket,      --                .endofpacket
			rf_source_data          => timer_0_s1_translator_avalon_universal_slave_0_agent_rf_source_data,             --                .data
			rdata_fifo_sink_ready   => timer_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready,       -- rdata_fifo_sink.ready
			rdata_fifo_sink_valid   => timer_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid,       --                .valid
			rdata_fifo_sink_data    => timer_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data,        --                .data
			rdata_fifo_src_ready    => timer_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready,       --  rdata_fifo_src.ready
			rdata_fifo_src_valid    => timer_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid,       --                .valid
			rdata_fifo_src_data     => timer_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data         --                .data
		);

	timer_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo : component Nios1_pio_LEDG_s1_translator_avalon_universal_slave_0_agent_rsp_fifo
		port map (
			clk               => clk_clk,                                                                         --       clk.clk
			reset             => rst_controller_reset_out_reset,                                                  -- clk_reset.reset
			in_data           => timer_0_s1_translator_avalon_universal_slave_0_agent_rf_source_data,             --        in.data
			in_valid          => timer_0_s1_translator_avalon_universal_slave_0_agent_rf_source_valid,            --          .valid
			in_ready          => timer_0_s1_translator_avalon_universal_slave_0_agent_rf_source_ready,            --          .ready
			in_startofpacket  => timer_0_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket,    --          .startofpacket
			in_endofpacket    => timer_0_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket,      --          .endofpacket
			out_data          => timer_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data,          --       out.data
			out_valid         => timer_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid,         --          .valid
			out_ready         => timer_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready,         --          .ready
			out_startofpacket => timer_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket, --          .startofpacket
			out_endofpacket   => timer_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket    --          .endofpacket
		);

	pio_rdydata_s1_translator_avalon_universal_slave_0_agent : component Nios1_pio_RdyData_s1_translator_avalon_universal_slave_0_agent
		port map (
			clk                     => clk_clk,                                                                             --             clk.clk
			reset                   => rst_controller_reset_out_reset,                                                      --       clk_reset.reset
			m0_address              => pio_rdydata_s1_translator_avalon_universal_slave_0_agent_m0_address,                 --              m0.address
			m0_burstcount           => pio_rdydata_s1_translator_avalon_universal_slave_0_agent_m0_burstcount,              --                .burstcount
			m0_byteenable           => pio_rdydata_s1_translator_avalon_universal_slave_0_agent_m0_byteenable,              --                .byteenable
			m0_debugaccess          => pio_rdydata_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess,             --                .debugaccess
			m0_lock                 => pio_rdydata_s1_translator_avalon_universal_slave_0_agent_m0_lock,                    --                .lock
			m0_readdata             => pio_rdydata_s1_translator_avalon_universal_slave_0_agent_m0_readdata,                --                .readdata
			m0_readdatavalid        => pio_rdydata_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid,           --                .readdatavalid
			m0_read                 => pio_rdydata_s1_translator_avalon_universal_slave_0_agent_m0_read,                    --                .read
			m0_waitrequest          => pio_rdydata_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest,             --                .waitrequest
			m0_writedata            => pio_rdydata_s1_translator_avalon_universal_slave_0_agent_m0_writedata,               --                .writedata
			m0_write                => pio_rdydata_s1_translator_avalon_universal_slave_0_agent_m0_write,                   --                .write
			rp_endofpacket          => pio_rdydata_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket,             --              rp.endofpacket
			rp_ready                => pio_rdydata_s1_translator_avalon_universal_slave_0_agent_rp_ready,                   --                .ready
			rp_valid                => pio_rdydata_s1_translator_avalon_universal_slave_0_agent_rp_valid,                   --                .valid
			rp_data                 => pio_rdydata_s1_translator_avalon_universal_slave_0_agent_rp_data,                    --                .data
			rp_startofpacket        => pio_rdydata_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket,           --                .startofpacket
			cp_ready                => cmd_xbar_demux_001_src12_ready,                                                      --              cp.ready
			cp_valid                => cmd_xbar_demux_001_src12_valid,                                                      --                .valid
			cp_data                 => cmd_xbar_demux_001_src12_data,                                                       --                .data
			cp_startofpacket        => cmd_xbar_demux_001_src12_startofpacket,                                              --                .startofpacket
			cp_endofpacket          => cmd_xbar_demux_001_src12_endofpacket,                                                --                .endofpacket
			cp_channel              => cmd_xbar_demux_001_src12_channel,                                                    --                .channel
			rf_sink_ready           => pio_rdydata_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready,         --         rf_sink.ready
			rf_sink_valid           => pio_rdydata_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid,         --                .valid
			rf_sink_startofpacket   => pio_rdydata_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket, --                .startofpacket
			rf_sink_endofpacket     => pio_rdydata_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket,   --                .endofpacket
			rf_sink_data            => pio_rdydata_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data,          --                .data
			rf_source_ready         => pio_rdydata_s1_translator_avalon_universal_slave_0_agent_rf_source_ready,            --       rf_source.ready
			rf_source_valid         => pio_rdydata_s1_translator_avalon_universal_slave_0_agent_rf_source_valid,            --                .valid
			rf_source_startofpacket => pio_rdydata_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket,    --                .startofpacket
			rf_source_endofpacket   => pio_rdydata_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket,      --                .endofpacket
			rf_source_data          => pio_rdydata_s1_translator_avalon_universal_slave_0_agent_rf_source_data,             --                .data
			rdata_fifo_sink_ready   => pio_rdydata_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready,       -- rdata_fifo_sink.ready
			rdata_fifo_sink_valid   => pio_rdydata_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid,       --                .valid
			rdata_fifo_sink_data    => pio_rdydata_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data,        --                .data
			rdata_fifo_src_ready    => pio_rdydata_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready,       --  rdata_fifo_src.ready
			rdata_fifo_src_valid    => pio_rdydata_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid,       --                .valid
			rdata_fifo_src_data     => pio_rdydata_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data         --                .data
		);

	pio_rdydata_s1_translator_avalon_universal_slave_0_agent_rsp_fifo : component Nios1_pio_LEDG_s1_translator_avalon_universal_slave_0_agent_rsp_fifo
		port map (
			clk               => clk_clk,                                                                             --       clk.clk
			reset             => rst_controller_reset_out_reset,                                                      -- clk_reset.reset
			in_data           => pio_rdydata_s1_translator_avalon_universal_slave_0_agent_rf_source_data,             --        in.data
			in_valid          => pio_rdydata_s1_translator_avalon_universal_slave_0_agent_rf_source_valid,            --          .valid
			in_ready          => pio_rdydata_s1_translator_avalon_universal_slave_0_agent_rf_source_ready,            --          .ready
			in_startofpacket  => pio_rdydata_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket,    --          .startofpacket
			in_endofpacket    => pio_rdydata_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket,      --          .endofpacket
			out_data          => pio_rdydata_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data,          --       out.data
			out_valid         => pio_rdydata_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid,         --          .valid
			out_ready         => pio_rdydata_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready,         --          .ready
			out_startofpacket => pio_rdydata_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket, --          .startofpacket
			out_endofpacket   => pio_rdydata_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket    --          .endofpacket
		);

	addr_router : component Nios1_addr_router
		port map (
			sink_ready         => nios2_qsys_instruction_master_translator_avalon_universal_master_0_agent_cp_ready,         --      sink.ready
			sink_valid         => nios2_qsys_instruction_master_translator_avalon_universal_master_0_agent_cp_valid,         --          .valid
			sink_data          => nios2_qsys_instruction_master_translator_avalon_universal_master_0_agent_cp_data,          --          .data
			sink_startofpacket => nios2_qsys_instruction_master_translator_avalon_universal_master_0_agent_cp_startofpacket, --          .startofpacket
			sink_endofpacket   => nios2_qsys_instruction_master_translator_avalon_universal_master_0_agent_cp_endofpacket,   --          .endofpacket
			clk                => clk_clk,                                                                                   --       clk.clk
			reset              => rst_controller_reset_out_reset,                                                            -- clk_reset.reset
			src_ready          => addr_router_src_ready,                                                                     --       src.ready
			src_valid          => addr_router_src_valid,                                                                     --          .valid
			src_data           => addr_router_src_data,                                                                      --          .data
			src_channel        => addr_router_src_channel,                                                                   --          .channel
			src_startofpacket  => addr_router_src_startofpacket,                                                             --          .startofpacket
			src_endofpacket    => addr_router_src_endofpacket                                                                --          .endofpacket
		);

	addr_router_001 : component Nios1_addr_router_001
		port map (
			sink_ready         => nios2_qsys_data_master_translator_avalon_universal_master_0_agent_cp_ready,         --      sink.ready
			sink_valid         => nios2_qsys_data_master_translator_avalon_universal_master_0_agent_cp_valid,         --          .valid
			sink_data          => nios2_qsys_data_master_translator_avalon_universal_master_0_agent_cp_data,          --          .data
			sink_startofpacket => nios2_qsys_data_master_translator_avalon_universal_master_0_agent_cp_startofpacket, --          .startofpacket
			sink_endofpacket   => nios2_qsys_data_master_translator_avalon_universal_master_0_agent_cp_endofpacket,   --          .endofpacket
			clk                => clk_clk,                                                                            --       clk.clk
			reset              => rst_controller_reset_out_reset,                                                     -- clk_reset.reset
			src_ready          => addr_router_001_src_ready,                                                          --       src.ready
			src_valid          => addr_router_001_src_valid,                                                          --          .valid
			src_data           => addr_router_001_src_data,                                                           --          .data
			src_channel        => addr_router_001_src_channel,                                                        --          .channel
			src_startofpacket  => addr_router_001_src_startofpacket,                                                  --          .startofpacket
			src_endofpacket    => addr_router_001_src_endofpacket                                                     --          .endofpacket
		);

	id_router : component Nios1_id_router
		port map (
			sink_ready         => nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_ready,         --      sink.ready
			sink_valid         => nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_valid,         --          .valid
			sink_data          => nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_data,          --          .data
			sink_startofpacket => nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_startofpacket, --          .startofpacket
			sink_endofpacket   => nios2_qsys_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_endofpacket,   --          .endofpacket
			clk                => clk_clk,                                                                                 --       clk.clk
			reset              => rst_controller_reset_out_reset,                                                          -- clk_reset.reset
			src_ready          => id_router_src_ready,                                                                     --       src.ready
			src_valid          => id_router_src_valid,                                                                     --          .valid
			src_data           => id_router_src_data,                                                                      --          .data
			src_channel        => id_router_src_channel,                                                                   --          .channel
			src_startofpacket  => id_router_src_startofpacket,                                                             --          .startofpacket
			src_endofpacket    => id_router_src_endofpacket                                                                --          .endofpacket
		);

	id_router_001 : component Nios1_id_router
		port map (
			sink_ready         => onchip_memory_s1_translator_avalon_universal_slave_0_agent_rp_ready,         --      sink.ready
			sink_valid         => onchip_memory_s1_translator_avalon_universal_slave_0_agent_rp_valid,         --          .valid
			sink_data          => onchip_memory_s1_translator_avalon_universal_slave_0_agent_rp_data,          --          .data
			sink_startofpacket => onchip_memory_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket, --          .startofpacket
			sink_endofpacket   => onchip_memory_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket,   --          .endofpacket
			clk                => clk_clk,                                                                     --       clk.clk
			reset              => rst_controller_reset_out_reset,                                              -- clk_reset.reset
			src_ready          => id_router_001_src_ready,                                                     --       src.ready
			src_valid          => id_router_001_src_valid,                                                     --          .valid
			src_data           => id_router_001_src_data,                                                      --          .data
			src_channel        => id_router_001_src_channel,                                                   --          .channel
			src_startofpacket  => id_router_001_src_startofpacket,                                             --          .startofpacket
			src_endofpacket    => id_router_001_src_endofpacket                                                --          .endofpacket
		);

	id_router_002 : component Nios1_id_router_002
		port map (
			sink_ready         => jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_ready,         --      sink.ready
			sink_valid         => jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_valid,         --          .valid
			sink_data          => jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_data,          --          .data
			sink_startofpacket => jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket, --          .startofpacket
			sink_endofpacket   => jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket,   --          .endofpacket
			clk                => clk_clk,                                                                                --       clk.clk
			reset              => rst_controller_reset_out_reset,                                                         -- clk_reset.reset
			src_ready          => id_router_002_src_ready,                                                                --       src.ready
			src_valid          => id_router_002_src_valid,                                                                --          .valid
			src_data           => id_router_002_src_data,                                                                 --          .data
			src_channel        => id_router_002_src_channel,                                                              --          .channel
			src_startofpacket  => id_router_002_src_startofpacket,                                                        --          .startofpacket
			src_endofpacket    => id_router_002_src_endofpacket                                                           --          .endofpacket
		);

	id_router_003 : component Nios1_id_router_002
		port map (
			sink_ready         => sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent_rp_ready,         --      sink.ready
			sink_valid         => sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent_rp_valid,         --          .valid
			sink_data          => sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent_rp_data,          --          .data
			sink_startofpacket => sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket, --          .startofpacket
			sink_endofpacket   => sysid_qsys_control_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket,   --          .endofpacket
			clk                => clk_clk,                                                                             --       clk.clk
			reset              => rst_controller_reset_out_reset,                                                      -- clk_reset.reset
			src_ready          => id_router_003_src_ready,                                                             --       src.ready
			src_valid          => id_router_003_src_valid,                                                             --          .valid
			src_data           => id_router_003_src_data,                                                              --          .data
			src_channel        => id_router_003_src_channel,                                                           --          .channel
			src_startofpacket  => id_router_003_src_startofpacket,                                                     --          .startofpacket
			src_endofpacket    => id_router_003_src_endofpacket                                                        --          .endofpacket
		);

	id_router_004 : component Nios1_id_router_002
		port map (
			sink_ready         => pio_ledg_s1_translator_avalon_universal_slave_0_agent_rp_ready,         --      sink.ready
			sink_valid         => pio_ledg_s1_translator_avalon_universal_slave_0_agent_rp_valid,         --          .valid
			sink_data          => pio_ledg_s1_translator_avalon_universal_slave_0_agent_rp_data,          --          .data
			sink_startofpacket => pio_ledg_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket, --          .startofpacket
			sink_endofpacket   => pio_ledg_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket,   --          .endofpacket
			clk                => clk_clk,                                                                --       clk.clk
			reset              => rst_controller_reset_out_reset,                                         -- clk_reset.reset
			src_ready          => id_router_004_src_ready,                                                --       src.ready
			src_valid          => id_router_004_src_valid,                                                --          .valid
			src_data           => id_router_004_src_data,                                                 --          .data
			src_channel        => id_router_004_src_channel,                                              --          .channel
			src_startofpacket  => id_router_004_src_startofpacket,                                        --          .startofpacket
			src_endofpacket    => id_router_004_src_endofpacket                                           --          .endofpacket
		);

	id_router_005 : component Nios1_id_router_002
		port map (
			sink_ready         => pio_ledr_s1_translator_avalon_universal_slave_0_agent_rp_ready,         --      sink.ready
			sink_valid         => pio_ledr_s1_translator_avalon_universal_slave_0_agent_rp_valid,         --          .valid
			sink_data          => pio_ledr_s1_translator_avalon_universal_slave_0_agent_rp_data,          --          .data
			sink_startofpacket => pio_ledr_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket, --          .startofpacket
			sink_endofpacket   => pio_ledr_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket,   --          .endofpacket
			clk                => clk_clk,                                                                --       clk.clk
			reset              => rst_controller_reset_out_reset,                                         -- clk_reset.reset
			src_ready          => id_router_005_src_ready,                                                --       src.ready
			src_valid          => id_router_005_src_valid,                                                --          .valid
			src_data           => id_router_005_src_data,                                                 --          .data
			src_channel        => id_router_005_src_channel,                                              --          .channel
			src_startofpacket  => id_router_005_src_startofpacket,                                        --          .startofpacket
			src_endofpacket    => id_router_005_src_endofpacket                                           --          .endofpacket
		);

	id_router_006 : component Nios1_id_router_002
		port map (
			sink_ready         => pio_sw_s1_translator_avalon_universal_slave_0_agent_rp_ready,         --      sink.ready
			sink_valid         => pio_sw_s1_translator_avalon_universal_slave_0_agent_rp_valid,         --          .valid
			sink_data          => pio_sw_s1_translator_avalon_universal_slave_0_agent_rp_data,          --          .data
			sink_startofpacket => pio_sw_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket, --          .startofpacket
			sink_endofpacket   => pio_sw_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket,   --          .endofpacket
			clk                => clk_clk,                                                              --       clk.clk
			reset              => rst_controller_reset_out_reset,                                       -- clk_reset.reset
			src_ready          => id_router_006_src_ready,                                              --       src.ready
			src_valid          => id_router_006_src_valid,                                              --          .valid
			src_data           => id_router_006_src_data,                                               --          .data
			src_channel        => id_router_006_src_channel,                                            --          .channel
			src_startofpacket  => id_router_006_src_startofpacket,                                      --          .startofpacket
			src_endofpacket    => id_router_006_src_endofpacket                                         --          .endofpacket
		);

	id_router_007 : component Nios1_id_router_002
		port map (
			sink_ready         => pio_button_s1_translator_avalon_universal_slave_0_agent_rp_ready,         --      sink.ready
			sink_valid         => pio_button_s1_translator_avalon_universal_slave_0_agent_rp_valid,         --          .valid
			sink_data          => pio_button_s1_translator_avalon_universal_slave_0_agent_rp_data,          --          .data
			sink_startofpacket => pio_button_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket, --          .startofpacket
			sink_endofpacket   => pio_button_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket,   --          .endofpacket
			clk                => clk_clk,                                                                  --       clk.clk
			reset              => rst_controller_reset_out_reset,                                           -- clk_reset.reset
			src_ready          => id_router_007_src_ready,                                                  --       src.ready
			src_valid          => id_router_007_src_valid,                                                  --          .valid
			src_data           => id_router_007_src_data,                                                   --          .data
			src_channel        => id_router_007_src_channel,                                                --          .channel
			src_startofpacket  => id_router_007_src_startofpacket,                                          --          .startofpacket
			src_endofpacket    => id_router_007_src_endofpacket                                             --          .endofpacket
		);

	id_router_008 : component Nios1_id_router_002
		port map (
			sink_ready         => lcd_control_slave_translator_avalon_universal_slave_0_agent_rp_ready,         --      sink.ready
			sink_valid         => lcd_control_slave_translator_avalon_universal_slave_0_agent_rp_valid,         --          .valid
			sink_data          => lcd_control_slave_translator_avalon_universal_slave_0_agent_rp_data,          --          .data
			sink_startofpacket => lcd_control_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket, --          .startofpacket
			sink_endofpacket   => lcd_control_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket,   --          .endofpacket
			clk                => clk_clk,                                                                      --       clk.clk
			reset              => rst_controller_reset_out_reset,                                               -- clk_reset.reset
			src_ready          => id_router_008_src_ready,                                                      --       src.ready
			src_valid          => id_router_008_src_valid,                                                      --          .valid
			src_data           => id_router_008_src_data,                                                       --          .data
			src_channel        => id_router_008_src_channel,                                                    --          .channel
			src_startofpacket  => id_router_008_src_startofpacket,                                              --          .startofpacket
			src_endofpacket    => id_router_008_src_endofpacket                                                 --          .endofpacket
		);

	id_router_009 : component Nios1_id_router_002
		port map (
			sink_ready         => uart_s1_translator_avalon_universal_slave_0_agent_rp_ready,         --      sink.ready
			sink_valid         => uart_s1_translator_avalon_universal_slave_0_agent_rp_valid,         --          .valid
			sink_data          => uart_s1_translator_avalon_universal_slave_0_agent_rp_data,          --          .data
			sink_startofpacket => uart_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket, --          .startofpacket
			sink_endofpacket   => uart_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket,   --          .endofpacket
			clk                => clk_clk,                                                            --       clk.clk
			reset              => rst_controller_reset_out_reset,                                     -- clk_reset.reset
			src_ready          => id_router_009_src_ready,                                            --       src.ready
			src_valid          => id_router_009_src_valid,                                            --          .valid
			src_data           => id_router_009_src_data,                                             --          .data
			src_channel        => id_router_009_src_channel,                                          --          .channel
			src_startofpacket  => id_router_009_src_startofpacket,                                    --          .startofpacket
			src_endofpacket    => id_router_009_src_endofpacket                                       --          .endofpacket
		);

	id_router_010 : component Nios1_id_router_002
		port map (
			sink_ready         => timer_0_s1_translator_avalon_universal_slave_0_agent_rp_ready,         --      sink.ready
			sink_valid         => timer_0_s1_translator_avalon_universal_slave_0_agent_rp_valid,         --          .valid
			sink_data          => timer_0_s1_translator_avalon_universal_slave_0_agent_rp_data,          --          .data
			sink_startofpacket => timer_0_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket, --          .startofpacket
			sink_endofpacket   => timer_0_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket,   --          .endofpacket
			clk                => clk_clk,                                                               --       clk.clk
			reset              => rst_controller_reset_out_reset,                                        -- clk_reset.reset
			src_ready          => id_router_010_src_ready,                                               --       src.ready
			src_valid          => id_router_010_src_valid,                                               --          .valid
			src_data           => id_router_010_src_data,                                                --          .data
			src_channel        => id_router_010_src_channel,                                             --          .channel
			src_startofpacket  => id_router_010_src_startofpacket,                                       --          .startofpacket
			src_endofpacket    => id_router_010_src_endofpacket                                          --          .endofpacket
		);

	id_router_011 : component Nios1_id_router_002
		port map (
			sink_ready         => pio_data_s1_translator_avalon_universal_slave_0_agent_rp_ready,         --      sink.ready
			sink_valid         => pio_data_s1_translator_avalon_universal_slave_0_agent_rp_valid,         --          .valid
			sink_data          => pio_data_s1_translator_avalon_universal_slave_0_agent_rp_data,          --          .data
			sink_startofpacket => pio_data_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket, --          .startofpacket
			sink_endofpacket   => pio_data_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket,   --          .endofpacket
			clk                => clk_clk,                                                                --       clk.clk
			reset              => rst_controller_reset_out_reset,                                         -- clk_reset.reset
			src_ready          => id_router_011_src_ready,                                                --       src.ready
			src_valid          => id_router_011_src_valid,                                                --          .valid
			src_data           => id_router_011_src_data,                                                 --          .data
			src_channel        => id_router_011_src_channel,                                              --          .channel
			src_startofpacket  => id_router_011_src_startofpacket,                                        --          .startofpacket
			src_endofpacket    => id_router_011_src_endofpacket                                           --          .endofpacket
		);

	id_router_012 : component Nios1_id_router_002
		port map (
			sink_ready         => pio_rdydata_s1_translator_avalon_universal_slave_0_agent_rp_ready,         --      sink.ready
			sink_valid         => pio_rdydata_s1_translator_avalon_universal_slave_0_agent_rp_valid,         --          .valid
			sink_data          => pio_rdydata_s1_translator_avalon_universal_slave_0_agent_rp_data,          --          .data
			sink_startofpacket => pio_rdydata_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket, --          .startofpacket
			sink_endofpacket   => pio_rdydata_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket,   --          .endofpacket
			clk                => clk_clk,                                                                   --       clk.clk
			reset              => rst_controller_reset_out_reset,                                            -- clk_reset.reset
			src_ready          => id_router_012_src_ready,                                                   --       src.ready
			src_valid          => id_router_012_src_valid,                                                   --          .valid
			src_data           => id_router_012_src_data,                                                    --          .data
			src_channel        => id_router_012_src_channel,                                                 --          .channel
			src_startofpacket  => id_router_012_src_startofpacket,                                           --          .startofpacket
			src_endofpacket    => id_router_012_src_endofpacket                                              --          .endofpacket
		);

	id_router_013 : component Nios1_id_router_002
		port map (
			sink_ready         => pio_dataread_s1_translator_avalon_universal_slave_0_agent_rp_ready,         --      sink.ready
			sink_valid         => pio_dataread_s1_translator_avalon_universal_slave_0_agent_rp_valid,         --          .valid
			sink_data          => pio_dataread_s1_translator_avalon_universal_slave_0_agent_rp_data,          --          .data
			sink_startofpacket => pio_dataread_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket, --          .startofpacket
			sink_endofpacket   => pio_dataread_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket,   --          .endofpacket
			clk                => clk_clk,                                                                    --       clk.clk
			reset              => rst_controller_reset_out_reset,                                             -- clk_reset.reset
			src_ready          => id_router_013_src_ready,                                                    --       src.ready
			src_valid          => id_router_013_src_valid,                                                    --          .valid
			src_data           => id_router_013_src_data,                                                     --          .data
			src_channel        => id_router_013_src_channel,                                                  --          .channel
			src_startofpacket  => id_router_013_src_startofpacket,                                            --          .startofpacket
			src_endofpacket    => id_router_013_src_endofpacket                                               --          .endofpacket
		);

	limiter : component Nios1_limiter
		port map (
			clk                    => clk_clk,                        --       clk.clk
			reset                  => rst_controller_reset_out_reset, -- clk_reset.reset
			cmd_sink_ready         => addr_router_src_ready,          --  cmd_sink.ready
			cmd_sink_valid         => addr_router_src_valid,          --          .valid
			cmd_sink_data          => addr_router_src_data,           --          .data
			cmd_sink_channel       => addr_router_src_channel,        --          .channel
			cmd_sink_startofpacket => addr_router_src_startofpacket,  --          .startofpacket
			cmd_sink_endofpacket   => addr_router_src_endofpacket,    --          .endofpacket
			cmd_src_ready          => limiter_cmd_src_ready,          --   cmd_src.ready
			cmd_src_data           => limiter_cmd_src_data,           --          .data
			cmd_src_channel        => limiter_cmd_src_channel,        --          .channel
			cmd_src_startofpacket  => limiter_cmd_src_startofpacket,  --          .startofpacket
			cmd_src_endofpacket    => limiter_cmd_src_endofpacket,    --          .endofpacket
			rsp_sink_ready         => rsp_xbar_mux_src_ready,         --  rsp_sink.ready
			rsp_sink_valid         => rsp_xbar_mux_src_valid,         --          .valid
			rsp_sink_channel       => rsp_xbar_mux_src_channel,       --          .channel
			rsp_sink_data          => rsp_xbar_mux_src_data,          --          .data
			rsp_sink_startofpacket => rsp_xbar_mux_src_startofpacket, --          .startofpacket
			rsp_sink_endofpacket   => rsp_xbar_mux_src_endofpacket,   --          .endofpacket
			rsp_src_ready          => limiter_rsp_src_ready,          --   rsp_src.ready
			rsp_src_valid          => limiter_rsp_src_valid,          --          .valid
			rsp_src_data           => limiter_rsp_src_data,           --          .data
			rsp_src_channel        => limiter_rsp_src_channel,        --          .channel
			rsp_src_startofpacket  => limiter_rsp_src_startofpacket,  --          .startofpacket
			rsp_src_endofpacket    => limiter_rsp_src_endofpacket,    --          .endofpacket
			cmd_src_valid          => limiter_cmd_valid_data          -- cmd_valid.data
		);

	limiter_001 : component Nios1_limiter
		port map (
			clk                    => clk_clk,                            --       clk.clk
			reset                  => rst_controller_reset_out_reset,     -- clk_reset.reset
			cmd_sink_ready         => addr_router_001_src_ready,          --  cmd_sink.ready
			cmd_sink_valid         => addr_router_001_src_valid,          --          .valid
			cmd_sink_data          => addr_router_001_src_data,           --          .data
			cmd_sink_channel       => addr_router_001_src_channel,        --          .channel
			cmd_sink_startofpacket => addr_router_001_src_startofpacket,  --          .startofpacket
			cmd_sink_endofpacket   => addr_router_001_src_endofpacket,    --          .endofpacket
			cmd_src_ready          => limiter_001_cmd_src_ready,          --   cmd_src.ready
			cmd_src_data           => limiter_001_cmd_src_data,           --          .data
			cmd_src_channel        => limiter_001_cmd_src_channel,        --          .channel
			cmd_src_startofpacket  => limiter_001_cmd_src_startofpacket,  --          .startofpacket
			cmd_src_endofpacket    => limiter_001_cmd_src_endofpacket,    --          .endofpacket
			rsp_sink_ready         => rsp_xbar_mux_001_src_ready,         --  rsp_sink.ready
			rsp_sink_valid         => rsp_xbar_mux_001_src_valid,         --          .valid
			rsp_sink_channel       => rsp_xbar_mux_001_src_channel,       --          .channel
			rsp_sink_data          => rsp_xbar_mux_001_src_data,          --          .data
			rsp_sink_startofpacket => rsp_xbar_mux_001_src_startofpacket, --          .startofpacket
			rsp_sink_endofpacket   => rsp_xbar_mux_001_src_endofpacket,   --          .endofpacket
			rsp_src_ready          => limiter_001_rsp_src_ready,          --   rsp_src.ready
			rsp_src_valid          => limiter_001_rsp_src_valid,          --          .valid
			rsp_src_data           => limiter_001_rsp_src_data,           --          .data
			rsp_src_channel        => limiter_001_rsp_src_channel,        --          .channel
			rsp_src_startofpacket  => limiter_001_rsp_src_startofpacket,  --          .startofpacket
			rsp_src_endofpacket    => limiter_001_rsp_src_endofpacket,    --          .endofpacket
			cmd_src_valid          => limiter_001_cmd_valid_data          -- cmd_valid.data
		);

	rst_controller : component Nios1_rst_controller
		port map (
			reset_in0 => reset_reset_n_ports_inv,        -- reset_in0.reset
			clk       => clk_clk,                        --       clk.clk
			reset_out => rst_controller_reset_out_reset  -- reset_out.reset
		);

	cmd_xbar_demux : component Nios1_cmd_xbar_demux
		port map (
			clk                => clk_clk,                           --        clk.clk
			reset              => rst_controller_reset_out_reset,    --  clk_reset.reset
			sink_ready         => limiter_cmd_src_ready,             --       sink.ready
			sink_channel       => limiter_cmd_src_channel,           --           .channel
			sink_data          => limiter_cmd_src_data,              --           .data
			sink_startofpacket => limiter_cmd_src_startofpacket,     --           .startofpacket
			sink_endofpacket   => limiter_cmd_src_endofpacket,       --           .endofpacket
			sink_valid         => limiter_cmd_valid_data,            -- sink_valid.data
			src0_ready         => cmd_xbar_demux_src0_ready,         --       src0.ready
			src0_valid         => cmd_xbar_demux_src0_valid,         --           .valid
			src0_data          => cmd_xbar_demux_src0_data,          --           .data
			src0_channel       => cmd_xbar_demux_src0_channel,       --           .channel
			src0_startofpacket => cmd_xbar_demux_src0_startofpacket, --           .startofpacket
			src0_endofpacket   => cmd_xbar_demux_src0_endofpacket,   --           .endofpacket
			src1_ready         => cmd_xbar_demux_src1_ready,         --       src1.ready
			src1_valid         => cmd_xbar_demux_src1_valid,         --           .valid
			src1_data          => cmd_xbar_demux_src1_data,          --           .data
			src1_channel       => cmd_xbar_demux_src1_channel,       --           .channel
			src1_startofpacket => cmd_xbar_demux_src1_startofpacket, --           .startofpacket
			src1_endofpacket   => cmd_xbar_demux_src1_endofpacket    --           .endofpacket
		);

	cmd_xbar_demux_001 : component Nios1_cmd_xbar_demux_001
		port map (
			clk                 => clk_clk,                                --        clk.clk
			reset               => rst_controller_reset_out_reset,         --  clk_reset.reset
			sink_ready          => limiter_001_cmd_src_ready,              --       sink.ready
			sink_channel        => limiter_001_cmd_src_channel,            --           .channel
			sink_data           => limiter_001_cmd_src_data,               --           .data
			sink_startofpacket  => limiter_001_cmd_src_startofpacket,      --           .startofpacket
			sink_endofpacket    => limiter_001_cmd_src_endofpacket,        --           .endofpacket
			sink_valid          => limiter_001_cmd_valid_data,             -- sink_valid.data
			src0_ready          => cmd_xbar_demux_001_src0_ready,          --       src0.ready
			src0_valid          => cmd_xbar_demux_001_src0_valid,          --           .valid
			src0_data           => cmd_xbar_demux_001_src0_data,           --           .data
			src0_channel        => cmd_xbar_demux_001_src0_channel,        --           .channel
			src0_startofpacket  => cmd_xbar_demux_001_src0_startofpacket,  --           .startofpacket
			src0_endofpacket    => cmd_xbar_demux_001_src0_endofpacket,    --           .endofpacket
			src1_ready          => cmd_xbar_demux_001_src1_ready,          --       src1.ready
			src1_valid          => cmd_xbar_demux_001_src1_valid,          --           .valid
			src1_data           => cmd_xbar_demux_001_src1_data,           --           .data
			src1_channel        => cmd_xbar_demux_001_src1_channel,        --           .channel
			src1_startofpacket  => cmd_xbar_demux_001_src1_startofpacket,  --           .startofpacket
			src1_endofpacket    => cmd_xbar_demux_001_src1_endofpacket,    --           .endofpacket
			src2_ready          => cmd_xbar_demux_001_src2_ready,          --       src2.ready
			src2_valid          => cmd_xbar_demux_001_src2_valid,          --           .valid
			src2_data           => cmd_xbar_demux_001_src2_data,           --           .data
			src2_channel        => cmd_xbar_demux_001_src2_channel,        --           .channel
			src2_startofpacket  => cmd_xbar_demux_001_src2_startofpacket,  --           .startofpacket
			src2_endofpacket    => cmd_xbar_demux_001_src2_endofpacket,    --           .endofpacket
			src3_ready          => cmd_xbar_demux_001_src3_ready,          --       src3.ready
			src3_valid          => cmd_xbar_demux_001_src3_valid,          --           .valid
			src3_data           => cmd_xbar_demux_001_src3_data,           --           .data
			src3_channel        => cmd_xbar_demux_001_src3_channel,        --           .channel
			src3_startofpacket  => cmd_xbar_demux_001_src3_startofpacket,  --           .startofpacket
			src3_endofpacket    => cmd_xbar_demux_001_src3_endofpacket,    --           .endofpacket
			src4_ready          => cmd_xbar_demux_001_src4_ready,          --       src4.ready
			src4_valid          => cmd_xbar_demux_001_src4_valid,          --           .valid
			src4_data           => cmd_xbar_demux_001_src4_data,           --           .data
			src4_channel        => cmd_xbar_demux_001_src4_channel,        --           .channel
			src4_startofpacket  => cmd_xbar_demux_001_src4_startofpacket,  --           .startofpacket
			src4_endofpacket    => cmd_xbar_demux_001_src4_endofpacket,    --           .endofpacket
			src5_ready          => cmd_xbar_demux_001_src5_ready,          --       src5.ready
			src5_valid          => cmd_xbar_demux_001_src5_valid,          --           .valid
			src5_data           => cmd_xbar_demux_001_src5_data,           --           .data
			src5_channel        => cmd_xbar_demux_001_src5_channel,        --           .channel
			src5_startofpacket  => cmd_xbar_demux_001_src5_startofpacket,  --           .startofpacket
			src5_endofpacket    => cmd_xbar_demux_001_src5_endofpacket,    --           .endofpacket
			src6_ready          => cmd_xbar_demux_001_src6_ready,          --       src6.ready
			src6_valid          => cmd_xbar_demux_001_src6_valid,          --           .valid
			src6_data           => cmd_xbar_demux_001_src6_data,           --           .data
			src6_channel        => cmd_xbar_demux_001_src6_channel,        --           .channel
			src6_startofpacket  => cmd_xbar_demux_001_src6_startofpacket,  --           .startofpacket
			src6_endofpacket    => cmd_xbar_demux_001_src6_endofpacket,    --           .endofpacket
			src7_ready          => cmd_xbar_demux_001_src7_ready,          --       src7.ready
			src7_valid          => cmd_xbar_demux_001_src7_valid,          --           .valid
			src7_data           => cmd_xbar_demux_001_src7_data,           --           .data
			src7_channel        => cmd_xbar_demux_001_src7_channel,        --           .channel
			src7_startofpacket  => cmd_xbar_demux_001_src7_startofpacket,  --           .startofpacket
			src7_endofpacket    => cmd_xbar_demux_001_src7_endofpacket,    --           .endofpacket
			src8_ready          => cmd_xbar_demux_001_src8_ready,          --       src8.ready
			src8_valid          => cmd_xbar_demux_001_src8_valid,          --           .valid
			src8_data           => cmd_xbar_demux_001_src8_data,           --           .data
			src8_channel        => cmd_xbar_demux_001_src8_channel,        --           .channel
			src8_startofpacket  => cmd_xbar_demux_001_src8_startofpacket,  --           .startofpacket
			src8_endofpacket    => cmd_xbar_demux_001_src8_endofpacket,    --           .endofpacket
			src9_ready          => cmd_xbar_demux_001_src9_ready,          --       src9.ready
			src9_valid          => cmd_xbar_demux_001_src9_valid,          --           .valid
			src9_data           => cmd_xbar_demux_001_src9_data,           --           .data
			src9_channel        => cmd_xbar_demux_001_src9_channel,        --           .channel
			src9_startofpacket  => cmd_xbar_demux_001_src9_startofpacket,  --           .startofpacket
			src9_endofpacket    => cmd_xbar_demux_001_src9_endofpacket,    --           .endofpacket
			src10_ready         => cmd_xbar_demux_001_src10_ready,         --      src10.ready
			src10_valid         => cmd_xbar_demux_001_src10_valid,         --           .valid
			src10_data          => cmd_xbar_demux_001_src10_data,          --           .data
			src10_channel       => cmd_xbar_demux_001_src10_channel,       --           .channel
			src10_startofpacket => cmd_xbar_demux_001_src10_startofpacket, --           .startofpacket
			src10_endofpacket   => cmd_xbar_demux_001_src10_endofpacket,   --           .endofpacket
			src11_ready         => cmd_xbar_demux_001_src11_ready,         --      src11.ready
			src11_valid         => cmd_xbar_demux_001_src11_valid,         --           .valid
			src11_data          => cmd_xbar_demux_001_src11_data,          --           .data
			src11_channel       => cmd_xbar_demux_001_src11_channel,       --           .channel
			src11_startofpacket => cmd_xbar_demux_001_src11_startofpacket, --           .startofpacket
			src11_endofpacket   => cmd_xbar_demux_001_src11_endofpacket,   --           .endofpacket
			src12_ready         => cmd_xbar_demux_001_src12_ready,         --      src12.ready
			src12_valid         => cmd_xbar_demux_001_src12_valid,         --           .valid
			src12_data          => cmd_xbar_demux_001_src12_data,          --           .data
			src12_channel       => cmd_xbar_demux_001_src12_channel,       --           .channel
			src12_startofpacket => cmd_xbar_demux_001_src12_startofpacket, --           .startofpacket
			src12_endofpacket   => cmd_xbar_demux_001_src12_endofpacket,   --           .endofpacket
			src13_ready         => cmd_xbar_demux_001_src13_ready,         --      src13.ready
			src13_valid         => cmd_xbar_demux_001_src13_valid,         --           .valid
			src13_data          => cmd_xbar_demux_001_src13_data,          --           .data
			src13_channel       => cmd_xbar_demux_001_src13_channel,       --           .channel
			src13_startofpacket => cmd_xbar_demux_001_src13_startofpacket, --           .startofpacket
			src13_endofpacket   => cmd_xbar_demux_001_src13_endofpacket    --           .endofpacket
		);

	cmd_xbar_mux : component Nios1_cmd_xbar_mux
		port map (
			clk                 => clk_clk,                               --       clk.clk
			reset               => rst_controller_reset_out_reset,        -- clk_reset.reset
			src_ready           => cmd_xbar_mux_src_ready,                --       src.ready
			src_valid           => cmd_xbar_mux_src_valid,                --          .valid
			src_data            => cmd_xbar_mux_src_data,                 --          .data
			src_channel         => cmd_xbar_mux_src_channel,              --          .channel
			src_startofpacket   => cmd_xbar_mux_src_startofpacket,        --          .startofpacket
			src_endofpacket     => cmd_xbar_mux_src_endofpacket,          --          .endofpacket
			sink0_ready         => cmd_xbar_demux_src0_ready,             --     sink0.ready
			sink0_valid         => cmd_xbar_demux_src0_valid,             --          .valid
			sink0_channel       => cmd_xbar_demux_src0_channel,           --          .channel
			sink0_data          => cmd_xbar_demux_src0_data,              --          .data
			sink0_startofpacket => cmd_xbar_demux_src0_startofpacket,     --          .startofpacket
			sink0_endofpacket   => cmd_xbar_demux_src0_endofpacket,       --          .endofpacket
			sink1_ready         => cmd_xbar_demux_001_src0_ready,         --     sink1.ready
			sink1_valid         => cmd_xbar_demux_001_src0_valid,         --          .valid
			sink1_channel       => cmd_xbar_demux_001_src0_channel,       --          .channel
			sink1_data          => cmd_xbar_demux_001_src0_data,          --          .data
			sink1_startofpacket => cmd_xbar_demux_001_src0_startofpacket, --          .startofpacket
			sink1_endofpacket   => cmd_xbar_demux_001_src0_endofpacket    --          .endofpacket
		);

	cmd_xbar_mux_001 : component Nios1_cmd_xbar_mux
		port map (
			clk                 => clk_clk,                               --       clk.clk
			reset               => rst_controller_reset_out_reset,        -- clk_reset.reset
			src_ready           => cmd_xbar_mux_001_src_ready,            --       src.ready
			src_valid           => cmd_xbar_mux_001_src_valid,            --          .valid
			src_data            => cmd_xbar_mux_001_src_data,             --          .data
			src_channel         => cmd_xbar_mux_001_src_channel,          --          .channel
			src_startofpacket   => cmd_xbar_mux_001_src_startofpacket,    --          .startofpacket
			src_endofpacket     => cmd_xbar_mux_001_src_endofpacket,      --          .endofpacket
			sink0_ready         => cmd_xbar_demux_src1_ready,             --     sink0.ready
			sink0_valid         => cmd_xbar_demux_src1_valid,             --          .valid
			sink0_channel       => cmd_xbar_demux_src1_channel,           --          .channel
			sink0_data          => cmd_xbar_demux_src1_data,              --          .data
			sink0_startofpacket => cmd_xbar_demux_src1_startofpacket,     --          .startofpacket
			sink0_endofpacket   => cmd_xbar_demux_src1_endofpacket,       --          .endofpacket
			sink1_ready         => cmd_xbar_demux_001_src1_ready,         --     sink1.ready
			sink1_valid         => cmd_xbar_demux_001_src1_valid,         --          .valid
			sink1_channel       => cmd_xbar_demux_001_src1_channel,       --          .channel
			sink1_data          => cmd_xbar_demux_001_src1_data,          --          .data
			sink1_startofpacket => cmd_xbar_demux_001_src1_startofpacket, --          .startofpacket
			sink1_endofpacket   => cmd_xbar_demux_001_src1_endofpacket    --          .endofpacket
		);

	rsp_xbar_demux : component Nios1_rsp_xbar_demux
		port map (
			clk                => clk_clk,                           --       clk.clk
			reset              => rst_controller_reset_out_reset,    -- clk_reset.reset
			sink_ready         => id_router_src_ready,               --      sink.ready
			sink_channel       => id_router_src_channel,             --          .channel
			sink_data          => id_router_src_data,                --          .data
			sink_startofpacket => id_router_src_startofpacket,       --          .startofpacket
			sink_endofpacket   => id_router_src_endofpacket,         --          .endofpacket
			sink_valid(0)      => id_router_src_valid,               --          .valid
			src0_ready         => rsp_xbar_demux_src0_ready,         --      src0.ready
			src0_valid         => rsp_xbar_demux_src0_valid,         --          .valid
			src0_data          => rsp_xbar_demux_src0_data,          --          .data
			src0_channel       => rsp_xbar_demux_src0_channel,       --          .channel
			src0_startofpacket => rsp_xbar_demux_src0_startofpacket, --          .startofpacket
			src0_endofpacket   => rsp_xbar_demux_src0_endofpacket,   --          .endofpacket
			src1_ready         => rsp_xbar_demux_src1_ready,         --      src1.ready
			src1_valid         => rsp_xbar_demux_src1_valid,         --          .valid
			src1_data          => rsp_xbar_demux_src1_data,          --          .data
			src1_channel       => rsp_xbar_demux_src1_channel,       --          .channel
			src1_startofpacket => rsp_xbar_demux_src1_startofpacket, --          .startofpacket
			src1_endofpacket   => rsp_xbar_demux_src1_endofpacket    --          .endofpacket
		);

	rsp_xbar_demux_001 : component Nios1_rsp_xbar_demux
		port map (
			clk                => clk_clk,                               --       clk.clk
			reset              => rst_controller_reset_out_reset,        -- clk_reset.reset
			sink_ready         => id_router_001_src_ready,               --      sink.ready
			sink_channel       => id_router_001_src_channel,             --          .channel
			sink_data          => id_router_001_src_data,                --          .data
			sink_startofpacket => id_router_001_src_startofpacket,       --          .startofpacket
			sink_endofpacket   => id_router_001_src_endofpacket,         --          .endofpacket
			sink_valid(0)      => id_router_001_src_valid,               --          .valid
			src0_ready         => rsp_xbar_demux_001_src0_ready,         --      src0.ready
			src0_valid         => rsp_xbar_demux_001_src0_valid,         --          .valid
			src0_data          => rsp_xbar_demux_001_src0_data,          --          .data
			src0_channel       => rsp_xbar_demux_001_src0_channel,       --          .channel
			src0_startofpacket => rsp_xbar_demux_001_src0_startofpacket, --          .startofpacket
			src0_endofpacket   => rsp_xbar_demux_001_src0_endofpacket,   --          .endofpacket
			src1_ready         => rsp_xbar_demux_001_src1_ready,         --      src1.ready
			src1_valid         => rsp_xbar_demux_001_src1_valid,         --          .valid
			src1_data          => rsp_xbar_demux_001_src1_data,          --          .data
			src1_channel       => rsp_xbar_demux_001_src1_channel,       --          .channel
			src1_startofpacket => rsp_xbar_demux_001_src1_startofpacket, --          .startofpacket
			src1_endofpacket   => rsp_xbar_demux_001_src1_endofpacket    --          .endofpacket
		);

	rsp_xbar_demux_002 : component Nios1_rsp_xbar_demux_002
		port map (
			clk                => clk_clk,                               --       clk.clk
			reset              => rst_controller_reset_out_reset,        -- clk_reset.reset
			sink_ready         => id_router_002_src_ready,               --      sink.ready
			sink_channel       => id_router_002_src_channel,             --          .channel
			sink_data          => id_router_002_src_data,                --          .data
			sink_startofpacket => id_router_002_src_startofpacket,       --          .startofpacket
			sink_endofpacket   => id_router_002_src_endofpacket,         --          .endofpacket
			sink_valid(0)      => id_router_002_src_valid,               --          .valid
			src0_ready         => rsp_xbar_demux_002_src0_ready,         --      src0.ready
			src0_valid         => rsp_xbar_demux_002_src0_valid,         --          .valid
			src0_data          => rsp_xbar_demux_002_src0_data,          --          .data
			src0_channel       => rsp_xbar_demux_002_src0_channel,       --          .channel
			src0_startofpacket => rsp_xbar_demux_002_src0_startofpacket, --          .startofpacket
			src0_endofpacket   => rsp_xbar_demux_002_src0_endofpacket    --          .endofpacket
		);

	rsp_xbar_demux_003 : component Nios1_rsp_xbar_demux_002
		port map (
			clk                => clk_clk,                               --       clk.clk
			reset              => rst_controller_reset_out_reset,        -- clk_reset.reset
			sink_ready         => id_router_003_src_ready,               --      sink.ready
			sink_channel       => id_router_003_src_channel,             --          .channel
			sink_data          => id_router_003_src_data,                --          .data
			sink_startofpacket => id_router_003_src_startofpacket,       --          .startofpacket
			sink_endofpacket   => id_router_003_src_endofpacket,         --          .endofpacket
			sink_valid(0)      => id_router_003_src_valid,               --          .valid
			src0_ready         => rsp_xbar_demux_003_src0_ready,         --      src0.ready
			src0_valid         => rsp_xbar_demux_003_src0_valid,         --          .valid
			src0_data          => rsp_xbar_demux_003_src0_data,          --          .data
			src0_channel       => rsp_xbar_demux_003_src0_channel,       --          .channel
			src0_startofpacket => rsp_xbar_demux_003_src0_startofpacket, --          .startofpacket
			src0_endofpacket   => rsp_xbar_demux_003_src0_endofpacket    --          .endofpacket
		);

	rsp_xbar_demux_004 : component Nios1_rsp_xbar_demux_002
		port map (
			clk                => clk_clk,                               --       clk.clk
			reset              => rst_controller_reset_out_reset,        -- clk_reset.reset
			sink_ready         => id_router_004_src_ready,               --      sink.ready
			sink_channel       => id_router_004_src_channel,             --          .channel
			sink_data          => id_router_004_src_data,                --          .data
			sink_startofpacket => id_router_004_src_startofpacket,       --          .startofpacket
			sink_endofpacket   => id_router_004_src_endofpacket,         --          .endofpacket
			sink_valid(0)      => id_router_004_src_valid,               --          .valid
			src0_ready         => rsp_xbar_demux_004_src0_ready,         --      src0.ready
			src0_valid         => rsp_xbar_demux_004_src0_valid,         --          .valid
			src0_data          => rsp_xbar_demux_004_src0_data,          --          .data
			src0_channel       => rsp_xbar_demux_004_src0_channel,       --          .channel
			src0_startofpacket => rsp_xbar_demux_004_src0_startofpacket, --          .startofpacket
			src0_endofpacket   => rsp_xbar_demux_004_src0_endofpacket    --          .endofpacket
		);

	rsp_xbar_demux_005 : component Nios1_rsp_xbar_demux_002
		port map (
			clk                => clk_clk,                               --       clk.clk
			reset              => rst_controller_reset_out_reset,        -- clk_reset.reset
			sink_ready         => id_router_005_src_ready,               --      sink.ready
			sink_channel       => id_router_005_src_channel,             --          .channel
			sink_data          => id_router_005_src_data,                --          .data
			sink_startofpacket => id_router_005_src_startofpacket,       --          .startofpacket
			sink_endofpacket   => id_router_005_src_endofpacket,         --          .endofpacket
			sink_valid(0)      => id_router_005_src_valid,               --          .valid
			src0_ready         => rsp_xbar_demux_005_src0_ready,         --      src0.ready
			src0_valid         => rsp_xbar_demux_005_src0_valid,         --          .valid
			src0_data          => rsp_xbar_demux_005_src0_data,          --          .data
			src0_channel       => rsp_xbar_demux_005_src0_channel,       --          .channel
			src0_startofpacket => rsp_xbar_demux_005_src0_startofpacket, --          .startofpacket
			src0_endofpacket   => rsp_xbar_demux_005_src0_endofpacket    --          .endofpacket
		);

	rsp_xbar_demux_006 : component Nios1_rsp_xbar_demux_002
		port map (
			clk                => clk_clk,                               --       clk.clk
			reset              => rst_controller_reset_out_reset,        -- clk_reset.reset
			sink_ready         => id_router_006_src_ready,               --      sink.ready
			sink_channel       => id_router_006_src_channel,             --          .channel
			sink_data          => id_router_006_src_data,                --          .data
			sink_startofpacket => id_router_006_src_startofpacket,       --          .startofpacket
			sink_endofpacket   => id_router_006_src_endofpacket,         --          .endofpacket
			sink_valid(0)      => id_router_006_src_valid,               --          .valid
			src0_ready         => rsp_xbar_demux_006_src0_ready,         --      src0.ready
			src0_valid         => rsp_xbar_demux_006_src0_valid,         --          .valid
			src0_data          => rsp_xbar_demux_006_src0_data,          --          .data
			src0_channel       => rsp_xbar_demux_006_src0_channel,       --          .channel
			src0_startofpacket => rsp_xbar_demux_006_src0_startofpacket, --          .startofpacket
			src0_endofpacket   => rsp_xbar_demux_006_src0_endofpacket    --          .endofpacket
		);

	rsp_xbar_demux_007 : component Nios1_rsp_xbar_demux_002
		port map (
			clk                => clk_clk,                               --       clk.clk
			reset              => rst_controller_reset_out_reset,        -- clk_reset.reset
			sink_ready         => id_router_007_src_ready,               --      sink.ready
			sink_channel       => id_router_007_src_channel,             --          .channel
			sink_data          => id_router_007_src_data,                --          .data
			sink_startofpacket => id_router_007_src_startofpacket,       --          .startofpacket
			sink_endofpacket   => id_router_007_src_endofpacket,         --          .endofpacket
			sink_valid(0)      => id_router_007_src_valid,               --          .valid
			src0_ready         => rsp_xbar_demux_007_src0_ready,         --      src0.ready
			src0_valid         => rsp_xbar_demux_007_src0_valid,         --          .valid
			src0_data          => rsp_xbar_demux_007_src0_data,          --          .data
			src0_channel       => rsp_xbar_demux_007_src0_channel,       --          .channel
			src0_startofpacket => rsp_xbar_demux_007_src0_startofpacket, --          .startofpacket
			src0_endofpacket   => rsp_xbar_demux_007_src0_endofpacket    --          .endofpacket
		);

	rsp_xbar_demux_008 : component Nios1_rsp_xbar_demux_002
		port map (
			clk                => clk_clk,                               --       clk.clk
			reset              => rst_controller_reset_out_reset,        -- clk_reset.reset
			sink_ready         => id_router_008_src_ready,               --      sink.ready
			sink_channel       => id_router_008_src_channel,             --          .channel
			sink_data          => id_router_008_src_data,                --          .data
			sink_startofpacket => id_router_008_src_startofpacket,       --          .startofpacket
			sink_endofpacket   => id_router_008_src_endofpacket,         --          .endofpacket
			sink_valid(0)      => id_router_008_src_valid,               --          .valid
			src0_ready         => rsp_xbar_demux_008_src0_ready,         --      src0.ready
			src0_valid         => rsp_xbar_demux_008_src0_valid,         --          .valid
			src0_data          => rsp_xbar_demux_008_src0_data,          --          .data
			src0_channel       => rsp_xbar_demux_008_src0_channel,       --          .channel
			src0_startofpacket => rsp_xbar_demux_008_src0_startofpacket, --          .startofpacket
			src0_endofpacket   => rsp_xbar_demux_008_src0_endofpacket    --          .endofpacket
		);

	rsp_xbar_demux_009 : component Nios1_rsp_xbar_demux_002
		port map (
			clk                => clk_clk,                               --       clk.clk
			reset              => rst_controller_reset_out_reset,        -- clk_reset.reset
			sink_ready         => id_router_009_src_ready,               --      sink.ready
			sink_channel       => id_router_009_src_channel,             --          .channel
			sink_data          => id_router_009_src_data,                --          .data
			sink_startofpacket => id_router_009_src_startofpacket,       --          .startofpacket
			sink_endofpacket   => id_router_009_src_endofpacket,         --          .endofpacket
			sink_valid(0)      => id_router_009_src_valid,               --          .valid
			src0_ready         => rsp_xbar_demux_009_src0_ready,         --      src0.ready
			src0_valid         => rsp_xbar_demux_009_src0_valid,         --          .valid
			src0_data          => rsp_xbar_demux_009_src0_data,          --          .data
			src0_channel       => rsp_xbar_demux_009_src0_channel,       --          .channel
			src0_startofpacket => rsp_xbar_demux_009_src0_startofpacket, --          .startofpacket
			src0_endofpacket   => rsp_xbar_demux_009_src0_endofpacket    --          .endofpacket
		);

	rsp_xbar_demux_010 : component Nios1_rsp_xbar_demux_002
		port map (
			clk                => clk_clk,                               --       clk.clk
			reset              => rst_controller_reset_out_reset,        -- clk_reset.reset
			sink_ready         => id_router_010_src_ready,               --      sink.ready
			sink_channel       => id_router_010_src_channel,             --          .channel
			sink_data          => id_router_010_src_data,                --          .data
			sink_startofpacket => id_router_010_src_startofpacket,       --          .startofpacket
			sink_endofpacket   => id_router_010_src_endofpacket,         --          .endofpacket
			sink_valid(0)      => id_router_010_src_valid,               --          .valid
			src0_ready         => rsp_xbar_demux_010_src0_ready,         --      src0.ready
			src0_valid         => rsp_xbar_demux_010_src0_valid,         --          .valid
			src0_data          => rsp_xbar_demux_010_src0_data,          --          .data
			src0_channel       => rsp_xbar_demux_010_src0_channel,       --          .channel
			src0_startofpacket => rsp_xbar_demux_010_src0_startofpacket, --          .startofpacket
			src0_endofpacket   => rsp_xbar_demux_010_src0_endofpacket    --          .endofpacket
		);

	rsp_xbar_demux_011 : component Nios1_rsp_xbar_demux_002
		port map (
			clk                => clk_clk,                               --       clk.clk
			reset              => rst_controller_reset_out_reset,        -- clk_reset.reset
			sink_ready         => id_router_011_src_ready,               --      sink.ready
			sink_channel       => id_router_011_src_channel,             --          .channel
			sink_data          => id_router_011_src_data,                --          .data
			sink_startofpacket => id_router_011_src_startofpacket,       --          .startofpacket
			sink_endofpacket   => id_router_011_src_endofpacket,         --          .endofpacket
			sink_valid(0)      => id_router_011_src_valid,               --          .valid
			src0_ready         => rsp_xbar_demux_011_src0_ready,         --      src0.ready
			src0_valid         => rsp_xbar_demux_011_src0_valid,         --          .valid
			src0_data          => rsp_xbar_demux_011_src0_data,          --          .data
			src0_channel       => rsp_xbar_demux_011_src0_channel,       --          .channel
			src0_startofpacket => rsp_xbar_demux_011_src0_startofpacket, --          .startofpacket
			src0_endofpacket   => rsp_xbar_demux_011_src0_endofpacket    --          .endofpacket
		);

	rsp_xbar_demux_012 : component Nios1_rsp_xbar_demux_002
		port map (
			clk                => clk_clk,                               --       clk.clk
			reset              => rst_controller_reset_out_reset,        -- clk_reset.reset
			sink_ready         => id_router_012_src_ready,               --      sink.ready
			sink_channel       => id_router_012_src_channel,             --          .channel
			sink_data          => id_router_012_src_data,                --          .data
			sink_startofpacket => id_router_012_src_startofpacket,       --          .startofpacket
			sink_endofpacket   => id_router_012_src_endofpacket,         --          .endofpacket
			sink_valid(0)      => id_router_012_src_valid,               --          .valid
			src0_ready         => rsp_xbar_demux_012_src0_ready,         --      src0.ready
			src0_valid         => rsp_xbar_demux_012_src0_valid,         --          .valid
			src0_data          => rsp_xbar_demux_012_src0_data,          --          .data
			src0_channel       => rsp_xbar_demux_012_src0_channel,       --          .channel
			src0_startofpacket => rsp_xbar_demux_012_src0_startofpacket, --          .startofpacket
			src0_endofpacket   => rsp_xbar_demux_012_src0_endofpacket    --          .endofpacket
		);

	rsp_xbar_demux_013 : component Nios1_rsp_xbar_demux_002
		port map (
			clk                => clk_clk,                               --       clk.clk
			reset              => rst_controller_reset_out_reset,        -- clk_reset.reset
			sink_ready         => id_router_013_src_ready,               --      sink.ready
			sink_channel       => id_router_013_src_channel,             --          .channel
			sink_data          => id_router_013_src_data,                --          .data
			sink_startofpacket => id_router_013_src_startofpacket,       --          .startofpacket
			sink_endofpacket   => id_router_013_src_endofpacket,         --          .endofpacket
			sink_valid(0)      => id_router_013_src_valid,               --          .valid
			src0_ready         => rsp_xbar_demux_013_src0_ready,         --      src0.ready
			src0_valid         => rsp_xbar_demux_013_src0_valid,         --          .valid
			src0_data          => rsp_xbar_demux_013_src0_data,          --          .data
			src0_channel       => rsp_xbar_demux_013_src0_channel,       --          .channel
			src0_startofpacket => rsp_xbar_demux_013_src0_startofpacket, --          .startofpacket
			src0_endofpacket   => rsp_xbar_demux_013_src0_endofpacket    --          .endofpacket
		);

	rsp_xbar_mux : component Nios1_rsp_xbar_mux
		port map (
			clk                 => clk_clk,                               --       clk.clk
			reset               => rst_controller_reset_out_reset,        -- clk_reset.reset
			src_ready           => rsp_xbar_mux_src_ready,                --       src.ready
			src_valid           => rsp_xbar_mux_src_valid,                --          .valid
			src_data            => rsp_xbar_mux_src_data,                 --          .data
			src_channel         => rsp_xbar_mux_src_channel,              --          .channel
			src_startofpacket   => rsp_xbar_mux_src_startofpacket,        --          .startofpacket
			src_endofpacket     => rsp_xbar_mux_src_endofpacket,          --          .endofpacket
			sink0_ready         => rsp_xbar_demux_src0_ready,             --     sink0.ready
			sink0_valid         => rsp_xbar_demux_src0_valid,             --          .valid
			sink0_channel       => rsp_xbar_demux_src0_channel,           --          .channel
			sink0_data          => rsp_xbar_demux_src0_data,              --          .data
			sink0_startofpacket => rsp_xbar_demux_src0_startofpacket,     --          .startofpacket
			sink0_endofpacket   => rsp_xbar_demux_src0_endofpacket,       --          .endofpacket
			sink1_ready         => rsp_xbar_demux_001_src0_ready,         --     sink1.ready
			sink1_valid         => rsp_xbar_demux_001_src0_valid,         --          .valid
			sink1_channel       => rsp_xbar_demux_001_src0_channel,       --          .channel
			sink1_data          => rsp_xbar_demux_001_src0_data,          --          .data
			sink1_startofpacket => rsp_xbar_demux_001_src0_startofpacket, --          .startofpacket
			sink1_endofpacket   => rsp_xbar_demux_001_src0_endofpacket    --          .endofpacket
		);

	rsp_xbar_mux_001 : component Nios1_rsp_xbar_mux_001
		port map (
			clk                  => clk_clk,                               --       clk.clk
			reset                => rst_controller_reset_out_reset,        -- clk_reset.reset
			src_ready            => rsp_xbar_mux_001_src_ready,            --       src.ready
			src_valid            => rsp_xbar_mux_001_src_valid,            --          .valid
			src_data             => rsp_xbar_mux_001_src_data,             --          .data
			src_channel          => rsp_xbar_mux_001_src_channel,          --          .channel
			src_startofpacket    => rsp_xbar_mux_001_src_startofpacket,    --          .startofpacket
			src_endofpacket      => rsp_xbar_mux_001_src_endofpacket,      --          .endofpacket
			sink0_ready          => rsp_xbar_demux_src1_ready,             --     sink0.ready
			sink0_valid          => rsp_xbar_demux_src1_valid,             --          .valid
			sink0_channel        => rsp_xbar_demux_src1_channel,           --          .channel
			sink0_data           => rsp_xbar_demux_src1_data,              --          .data
			sink0_startofpacket  => rsp_xbar_demux_src1_startofpacket,     --          .startofpacket
			sink0_endofpacket    => rsp_xbar_demux_src1_endofpacket,       --          .endofpacket
			sink1_ready          => rsp_xbar_demux_001_src1_ready,         --     sink1.ready
			sink1_valid          => rsp_xbar_demux_001_src1_valid,         --          .valid
			sink1_channel        => rsp_xbar_demux_001_src1_channel,       --          .channel
			sink1_data           => rsp_xbar_demux_001_src1_data,          --          .data
			sink1_startofpacket  => rsp_xbar_demux_001_src1_startofpacket, --          .startofpacket
			sink1_endofpacket    => rsp_xbar_demux_001_src1_endofpacket,   --          .endofpacket
			sink2_ready          => rsp_xbar_demux_002_src0_ready,         --     sink2.ready
			sink2_valid          => rsp_xbar_demux_002_src0_valid,         --          .valid
			sink2_channel        => rsp_xbar_demux_002_src0_channel,       --          .channel
			sink2_data           => rsp_xbar_demux_002_src0_data,          --          .data
			sink2_startofpacket  => rsp_xbar_demux_002_src0_startofpacket, --          .startofpacket
			sink2_endofpacket    => rsp_xbar_demux_002_src0_endofpacket,   --          .endofpacket
			sink3_ready          => rsp_xbar_demux_003_src0_ready,         --     sink3.ready
			sink3_valid          => rsp_xbar_demux_003_src0_valid,         --          .valid
			sink3_channel        => rsp_xbar_demux_003_src0_channel,       --          .channel
			sink3_data           => rsp_xbar_demux_003_src0_data,          --          .data
			sink3_startofpacket  => rsp_xbar_demux_003_src0_startofpacket, --          .startofpacket
			sink3_endofpacket    => rsp_xbar_demux_003_src0_endofpacket,   --          .endofpacket
			sink4_ready          => rsp_xbar_demux_004_src0_ready,         --     sink4.ready
			sink4_valid          => rsp_xbar_demux_004_src0_valid,         --          .valid
			sink4_channel        => rsp_xbar_demux_004_src0_channel,       --          .channel
			sink4_data           => rsp_xbar_demux_004_src0_data,          --          .data
			sink4_startofpacket  => rsp_xbar_demux_004_src0_startofpacket, --          .startofpacket
			sink4_endofpacket    => rsp_xbar_demux_004_src0_endofpacket,   --          .endofpacket
			sink5_ready          => rsp_xbar_demux_005_src0_ready,         --     sink5.ready
			sink5_valid          => rsp_xbar_demux_005_src0_valid,         --          .valid
			sink5_channel        => rsp_xbar_demux_005_src0_channel,       --          .channel
			sink5_data           => rsp_xbar_demux_005_src0_data,          --          .data
			sink5_startofpacket  => rsp_xbar_demux_005_src0_startofpacket, --          .startofpacket
			sink5_endofpacket    => rsp_xbar_demux_005_src0_endofpacket,   --          .endofpacket
			sink6_ready          => rsp_xbar_demux_006_src0_ready,         --     sink6.ready
			sink6_valid          => rsp_xbar_demux_006_src0_valid,         --          .valid
			sink6_channel        => rsp_xbar_demux_006_src0_channel,       --          .channel
			sink6_data           => rsp_xbar_demux_006_src0_data,          --          .data
			sink6_startofpacket  => rsp_xbar_demux_006_src0_startofpacket, --          .startofpacket
			sink6_endofpacket    => rsp_xbar_demux_006_src0_endofpacket,   --          .endofpacket
			sink7_ready          => rsp_xbar_demux_007_src0_ready,         --     sink7.ready
			sink7_valid          => rsp_xbar_demux_007_src0_valid,         --          .valid
			sink7_channel        => rsp_xbar_demux_007_src0_channel,       --          .channel
			sink7_data           => rsp_xbar_demux_007_src0_data,          --          .data
			sink7_startofpacket  => rsp_xbar_demux_007_src0_startofpacket, --          .startofpacket
			sink7_endofpacket    => rsp_xbar_demux_007_src0_endofpacket,   --          .endofpacket
			sink8_ready          => rsp_xbar_demux_008_src0_ready,         --     sink8.ready
			sink8_valid          => rsp_xbar_demux_008_src0_valid,         --          .valid
			sink8_channel        => rsp_xbar_demux_008_src0_channel,       --          .channel
			sink8_data           => rsp_xbar_demux_008_src0_data,          --          .data
			sink8_startofpacket  => rsp_xbar_demux_008_src0_startofpacket, --          .startofpacket
			sink8_endofpacket    => rsp_xbar_demux_008_src0_endofpacket,   --          .endofpacket
			sink9_ready          => rsp_xbar_demux_009_src0_ready,         --     sink9.ready
			sink9_valid          => rsp_xbar_demux_009_src0_valid,         --          .valid
			sink9_channel        => rsp_xbar_demux_009_src0_channel,       --          .channel
			sink9_data           => rsp_xbar_demux_009_src0_data,          --          .data
			sink9_startofpacket  => rsp_xbar_demux_009_src0_startofpacket, --          .startofpacket
			sink9_endofpacket    => rsp_xbar_demux_009_src0_endofpacket,   --          .endofpacket
			sink10_ready         => rsp_xbar_demux_010_src0_ready,         --    sink10.ready
			sink10_valid         => rsp_xbar_demux_010_src0_valid,         --          .valid
			sink10_channel       => rsp_xbar_demux_010_src0_channel,       --          .channel
			sink10_data          => rsp_xbar_demux_010_src0_data,          --          .data
			sink10_startofpacket => rsp_xbar_demux_010_src0_startofpacket, --          .startofpacket
			sink10_endofpacket   => rsp_xbar_demux_010_src0_endofpacket,   --          .endofpacket
			sink11_ready         => rsp_xbar_demux_011_src0_ready,         --    sink11.ready
			sink11_valid         => rsp_xbar_demux_011_src0_valid,         --          .valid
			sink11_channel       => rsp_xbar_demux_011_src0_channel,       --          .channel
			sink11_data          => rsp_xbar_demux_011_src0_data,          --          .data
			sink11_startofpacket => rsp_xbar_demux_011_src0_startofpacket, --          .startofpacket
			sink11_endofpacket   => rsp_xbar_demux_011_src0_endofpacket,   --          .endofpacket
			sink12_ready         => rsp_xbar_demux_012_src0_ready,         --    sink12.ready
			sink12_valid         => rsp_xbar_demux_012_src0_valid,         --          .valid
			sink12_channel       => rsp_xbar_demux_012_src0_channel,       --          .channel
			sink12_data          => rsp_xbar_demux_012_src0_data,          --          .data
			sink12_startofpacket => rsp_xbar_demux_012_src0_startofpacket, --          .startofpacket
			sink12_endofpacket   => rsp_xbar_demux_012_src0_endofpacket,   --          .endofpacket
			sink13_ready         => rsp_xbar_demux_013_src0_ready,         --    sink13.ready
			sink13_valid         => rsp_xbar_demux_013_src0_valid,         --          .valid
			sink13_channel       => rsp_xbar_demux_013_src0_channel,       --          .channel
			sink13_data          => rsp_xbar_demux_013_src0_data,          --          .data
			sink13_startofpacket => rsp_xbar_demux_013_src0_startofpacket, --          .startofpacket
			sink13_endofpacket   => rsp_xbar_demux_013_src0_endofpacket    --          .endofpacket
		);

	irq_mapper : component Nios1_irq_mapper
		port map (
			clk           => clk_clk,                        --       clk.clk
			reset         => rst_controller_reset_out_reset, -- clk_reset.reset
			receiver0_irq => irq_mapper_receiver0_irq,       -- receiver0.irq
			receiver1_irq => irq_mapper_receiver1_irq,       -- receiver1.irq
			receiver2_irq => irq_mapper_receiver2_irq,       -- receiver2.irq
			receiver3_irq => irq_mapper_receiver3_irq,       -- receiver3.irq
			receiver4_irq => irq_mapper_receiver4_irq,       -- receiver4.irq
			sender_irq    => nios2_qsys_d_irq_irq            --    sender.irq
		);

	reset_reset_n_ports_inv <= not reset_reset_n;

	jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_write_ports_inv <= not jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_write;

	jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_read_ports_inv <= not jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_read;

	pio_ledg_s1_translator_avalon_anti_slave_0_write_ports_inv <= not pio_ledg_s1_translator_avalon_anti_slave_0_write;

	pio_ledr_s1_translator_avalon_anti_slave_0_write_ports_inv <= not pio_ledr_s1_translator_avalon_anti_slave_0_write;

	pio_button_s1_translator_avalon_anti_slave_0_write_ports_inv <= not pio_button_s1_translator_avalon_anti_slave_0_write;

	uart_s1_translator_avalon_anti_slave_0_write_ports_inv <= not uart_s1_translator_avalon_anti_slave_0_write;

	uart_s1_translator_avalon_anti_slave_0_read_ports_inv <= not uart_s1_translator_avalon_anti_slave_0_read;

	timer_0_s1_translator_avalon_anti_slave_0_write_ports_inv <= not timer_0_s1_translator_avalon_anti_slave_0_write;

	pio_rdydata_s1_translator_avalon_anti_slave_0_write_ports_inv <= not pio_rdydata_s1_translator_avalon_anti_slave_0_write;

	pio_dataread_s1_translator_avalon_anti_slave_0_write_ports_inv <= not pio_dataread_s1_translator_avalon_anti_slave_0_write;

	rst_controller_reset_out_reset_ports_inv <= not rst_controller_reset_out_reset;

end architecture rtl; -- of Nios1
